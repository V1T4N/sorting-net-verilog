module sort_pipe(
     input clk,
     input  [7:0]x_0, x_1, x_2, x_3, x_4, x_5, x_6, x_7, x_8, x_9, x_10, x_11, x_12, x_13, x_14, x_15, x_16, x_17, x_18, x_19, x_20, x_21, x_22, x_23, x_24, x_25, x_26, x_27, x_28, x_29, x_30, x_31, x_32, x_33, x_34, x_35, x_36, x_37, x_38, x_39, x_40, x_41, x_42, x_43, x_44, x_45, x_46, x_47, x_48, 
     output [7:0] median
);
reg[7:0] r0 [48:0];
reg[7:0] r1 [48:0];
reg[7:0] r2 [48:0];
reg[7:0] r3 [48:0];
reg[7:0] r4 [48:0];
reg[7:0] r5 [48:0];
reg[7:0] r6 [48:0];
reg[7:0] r7 [48:0];
reg[7:0] r8 [48:0];
reg[7:0] r9 [48:0];
reg[7:0] r10 [48:0];
reg[7:0] r11 [48:0];
reg[7:0] r12 [48:0];
reg[7:0] r13 [48:0];
reg[7:0] r14 [48:0];
reg[7:0] r15 [48:0];
reg[7:0] r16 [48:0];
reg[7:0] r17 [48:0];
reg[7:0] r18 [48:0];
reg[7:0] r19 [48:0];
reg[7:0] r20 [48:0];

//-------dec layer:0----------
wire [7:0] cmp0_out0;
wire [7:0] cmp0_out1;
reg [7:0] cmp0_in0;
reg [7:0] cmp0_in1;

wire [7:0] cmp1_out0;
wire [7:0] cmp1_out1;
reg [7:0] cmp1_in0;
reg [7:0] cmp1_in1;

wire [7:0] cmp2_out0;
wire [7:0] cmp2_out1;
reg [7:0] cmp2_in0;
reg [7:0] cmp2_in1;

wire [7:0] cmp3_out0;
wire [7:0] cmp3_out1;
reg [7:0] cmp3_in0;
reg [7:0] cmp3_in1;

wire [7:0] cmp4_out0;
wire [7:0] cmp4_out1;
reg [7:0] cmp4_in0;
reg [7:0] cmp4_in1;

wire [7:0] cmp5_out0;
wire [7:0] cmp5_out1;
reg [7:0] cmp5_in0;
reg [7:0] cmp5_in1;

wire [7:0] cmp6_out0;
wire [7:0] cmp6_out1;
reg [7:0] cmp6_in0;
reg [7:0] cmp6_in1;

wire [7:0] cmp7_out0;
wire [7:0] cmp7_out1;
reg [7:0] cmp7_in0;
reg [7:0] cmp7_in1;

wire [7:0] cmp8_out0;
wire [7:0] cmp8_out1;
reg [7:0] cmp8_in0;
reg [7:0] cmp8_in1;

wire [7:0] cmp9_out0;
wire [7:0] cmp9_out1;
reg [7:0] cmp9_in0;
reg [7:0] cmp9_in1;

wire [7:0] cmp10_out0;
wire [7:0] cmp10_out1;
reg [7:0] cmp10_in0;
reg [7:0] cmp10_in1;

wire [7:0] cmp11_out0;
wire [7:0] cmp11_out1;
reg [7:0] cmp11_in0;
reg [7:0] cmp11_in1;

wire [7:0] cmp12_out0;
wire [7:0] cmp12_out1;
reg [7:0] cmp12_in0;
reg [7:0] cmp12_in1;

wire [7:0] cmp13_out0;
wire [7:0] cmp13_out1;
reg [7:0] cmp13_in0;
reg [7:0] cmp13_in1;

wire [7:0] cmp14_out0;
wire [7:0] cmp14_out1;
reg [7:0] cmp14_in0;
reg [7:0] cmp14_in1;

wire [7:0] cmp15_out0;
wire [7:0] cmp15_out1;
reg [7:0] cmp15_in0;
reg [7:0] cmp15_in1;

wire [7:0] cmp16_out0;
wire [7:0] cmp16_out1;
reg [7:0] cmp16_in0;
reg [7:0] cmp16_in1;

//-------dec layer:1----------
wire [7:0] cmp17_out0;
wire [7:0] cmp17_out1;
reg [7:0] cmp17_in0;
reg [7:0] cmp17_in1;

wire [7:0] cmp18_out0;
wire [7:0] cmp18_out1;
reg [7:0] cmp18_in0;
reg [7:0] cmp18_in1;

wire [7:0] cmp19_out0;
wire [7:0] cmp19_out1;
reg [7:0] cmp19_in0;
reg [7:0] cmp19_in1;

wire [7:0] cmp20_out0;
wire [7:0] cmp20_out1;
reg [7:0] cmp20_in0;
reg [7:0] cmp20_in1;

wire [7:0] cmp21_out0;
wire [7:0] cmp21_out1;
reg [7:0] cmp21_in0;
reg [7:0] cmp21_in1;

wire [7:0] cmp22_out0;
wire [7:0] cmp22_out1;
reg [7:0] cmp22_in0;
reg [7:0] cmp22_in1;

wire [7:0] cmp23_out0;
wire [7:0] cmp23_out1;
reg [7:0] cmp23_in0;
reg [7:0] cmp23_in1;

wire [7:0] cmp24_out0;
wire [7:0] cmp24_out1;
reg [7:0] cmp24_in0;
reg [7:0] cmp24_in1;

wire [7:0] cmp25_out0;
wire [7:0] cmp25_out1;
reg [7:0] cmp25_in0;
reg [7:0] cmp25_in1;

wire [7:0] cmp26_out0;
wire [7:0] cmp26_out1;
reg [7:0] cmp26_in0;
reg [7:0] cmp26_in1;

wire [7:0] cmp27_out0;
wire [7:0] cmp27_out1;
reg [7:0] cmp27_in0;
reg [7:0] cmp27_in1;

wire [7:0] cmp28_out0;
wire [7:0] cmp28_out1;
reg [7:0] cmp28_in0;
reg [7:0] cmp28_in1;

wire [7:0] cmp29_out0;
wire [7:0] cmp29_out1;
reg [7:0] cmp29_in0;
reg [7:0] cmp29_in1;

wire [7:0] cmp30_out0;
wire [7:0] cmp30_out1;
reg [7:0] cmp30_in0;
reg [7:0] cmp30_in1;

wire [7:0] cmp31_out0;
wire [7:0] cmp31_out1;
reg [7:0] cmp31_in0;
reg [7:0] cmp31_in1;

wire [7:0] cmp32_out0;
wire [7:0] cmp32_out1;
reg [7:0] cmp32_in0;
reg [7:0] cmp32_in1;

wire [7:0] cmp33_out0;
wire [7:0] cmp33_out1;
reg [7:0] cmp33_in0;
reg [7:0] cmp33_in1;

//-------dec layer:2----------
wire [7:0] cmp34_out0;
wire [7:0] cmp34_out1;
reg [7:0] cmp34_in0;
reg [7:0] cmp34_in1;

wire [7:0] cmp35_out0;
wire [7:0] cmp35_out1;
reg [7:0] cmp35_in0;
reg [7:0] cmp35_in1;

wire [7:0] cmp36_out0;
wire [7:0] cmp36_out1;
reg [7:0] cmp36_in0;
reg [7:0] cmp36_in1;

wire [7:0] cmp37_out0;
wire [7:0] cmp37_out1;
reg [7:0] cmp37_in0;
reg [7:0] cmp37_in1;

wire [7:0] cmp38_out0;
wire [7:0] cmp38_out1;
reg [7:0] cmp38_in0;
reg [7:0] cmp38_in1;

wire [7:0] cmp39_out0;
wire [7:0] cmp39_out1;
reg [7:0] cmp39_in0;
reg [7:0] cmp39_in1;

wire [7:0] cmp40_out0;
wire [7:0] cmp40_out1;
reg [7:0] cmp40_in0;
reg [7:0] cmp40_in1;

wire [7:0] cmp41_out0;
wire [7:0] cmp41_out1;
reg [7:0] cmp41_in0;
reg [7:0] cmp41_in1;

wire [7:0] cmp42_out0;
wire [7:0] cmp42_out1;
reg [7:0] cmp42_in0;
reg [7:0] cmp42_in1;

wire [7:0] cmp43_out0;
wire [7:0] cmp43_out1;
reg [7:0] cmp43_in0;
reg [7:0] cmp43_in1;

wire [7:0] cmp44_out0;
wire [7:0] cmp44_out1;
reg [7:0] cmp44_in0;
reg [7:0] cmp44_in1;

wire [7:0] cmp45_out0;
wire [7:0] cmp45_out1;
reg [7:0] cmp45_in0;
reg [7:0] cmp45_in1;

wire [7:0] cmp46_out0;
wire [7:0] cmp46_out1;
reg [7:0] cmp46_in0;
reg [7:0] cmp46_in1;

wire [7:0] cmp47_out0;
wire [7:0] cmp47_out1;
reg [7:0] cmp47_in0;
reg [7:0] cmp47_in1;

wire [7:0] cmp48_out0;
wire [7:0] cmp48_out1;
reg [7:0] cmp48_in0;
reg [7:0] cmp48_in1;

wire [7:0] cmp49_out0;
wire [7:0] cmp49_out1;
reg [7:0] cmp49_in0;
reg [7:0] cmp49_in1;

wire [7:0] cmp50_out0;
wire [7:0] cmp50_out1;
reg [7:0] cmp50_in0;
reg [7:0] cmp50_in1;

wire [7:0] cmp51_out0;
wire [7:0] cmp51_out1;
reg [7:0] cmp51_in0;
reg [7:0] cmp51_in1;

wire [7:0] cmp52_out0;
wire [7:0] cmp52_out1;
reg [7:0] cmp52_in0;
reg [7:0] cmp52_in1;

wire [7:0] cmp53_out0;
wire [7:0] cmp53_out1;
reg [7:0] cmp53_in0;
reg [7:0] cmp53_in1;

wire [7:0] cmp54_out0;
wire [7:0] cmp54_out1;
reg [7:0] cmp54_in0;
reg [7:0] cmp54_in1;

wire [7:0] cmp55_out0;
wire [7:0] cmp55_out1;
reg [7:0] cmp55_in0;
reg [7:0] cmp55_in1;

wire [7:0] cmp56_out0;
wire [7:0] cmp56_out1;
reg [7:0] cmp56_in0;
reg [7:0] cmp56_in1;

wire [7:0] cmp57_out0;
wire [7:0] cmp57_out1;
reg [7:0] cmp57_in0;
reg [7:0] cmp57_in1;

//-------dec layer:3----------
wire [7:0] cmp58_out0;
wire [7:0] cmp58_out1;
reg [7:0] cmp58_in0;
reg [7:0] cmp58_in1;

wire [7:0] cmp59_out0;
wire [7:0] cmp59_out1;
reg [7:0] cmp59_in0;
reg [7:0] cmp59_in1;

wire [7:0] cmp60_out0;
wire [7:0] cmp60_out1;
reg [7:0] cmp60_in0;
reg [7:0] cmp60_in1;

wire [7:0] cmp61_out0;
wire [7:0] cmp61_out1;
reg [7:0] cmp61_in0;
reg [7:0] cmp61_in1;

wire [7:0] cmp62_out0;
wire [7:0] cmp62_out1;
reg [7:0] cmp62_in0;
reg [7:0] cmp62_in1;

wire [7:0] cmp63_out0;
wire [7:0] cmp63_out1;
reg [7:0] cmp63_in0;
reg [7:0] cmp63_in1;

wire [7:0] cmp64_out0;
wire [7:0] cmp64_out1;
reg [7:0] cmp64_in0;
reg [7:0] cmp64_in1;

wire [7:0] cmp65_out0;
wire [7:0] cmp65_out1;
reg [7:0] cmp65_in0;
reg [7:0] cmp65_in1;

wire [7:0] cmp66_out0;
wire [7:0] cmp66_out1;
reg [7:0] cmp66_in0;
reg [7:0] cmp66_in1;

wire [7:0] cmp67_out0;
wire [7:0] cmp67_out1;
reg [7:0] cmp67_in0;
reg [7:0] cmp67_in1;

wire [7:0] cmp68_out0;
wire [7:0] cmp68_out1;
reg [7:0] cmp68_in0;
reg [7:0] cmp68_in1;

wire [7:0] cmp69_out0;
wire [7:0] cmp69_out1;
reg [7:0] cmp69_in0;
reg [7:0] cmp69_in1;

wire [7:0] cmp70_out0;
wire [7:0] cmp70_out1;
reg [7:0] cmp70_in0;
reg [7:0] cmp70_in1;

wire [7:0] cmp71_out0;
wire [7:0] cmp71_out1;
reg [7:0] cmp71_in0;
reg [7:0] cmp71_in1;

wire [7:0] cmp72_out0;
wire [7:0] cmp72_out1;
reg [7:0] cmp72_in0;
reg [7:0] cmp72_in1;

wire [7:0] cmp73_out0;
wire [7:0] cmp73_out1;
reg [7:0] cmp73_in0;
reg [7:0] cmp73_in1;

//-------dec layer:4----------
wire [7:0] cmp74_out0;
wire [7:0] cmp74_out1;
reg [7:0] cmp74_in0;
reg [7:0] cmp74_in1;

wire [7:0] cmp75_out0;
wire [7:0] cmp75_out1;
reg [7:0] cmp75_in0;
reg [7:0] cmp75_in1;

wire [7:0] cmp76_out0;
wire [7:0] cmp76_out1;
reg [7:0] cmp76_in0;
reg [7:0] cmp76_in1;

wire [7:0] cmp77_out0;
wire [7:0] cmp77_out1;
reg [7:0] cmp77_in0;
reg [7:0] cmp77_in1;

wire [7:0] cmp78_out0;
wire [7:0] cmp78_out1;
reg [7:0] cmp78_in0;
reg [7:0] cmp78_in1;

wire [7:0] cmp79_out0;
wire [7:0] cmp79_out1;
reg [7:0] cmp79_in0;
reg [7:0] cmp79_in1;

wire [7:0] cmp80_out0;
wire [7:0] cmp80_out1;
reg [7:0] cmp80_in0;
reg [7:0] cmp80_in1;

wire [7:0] cmp81_out0;
wire [7:0] cmp81_out1;
reg [7:0] cmp81_in0;
reg [7:0] cmp81_in1;

wire [7:0] cmp82_out0;
wire [7:0] cmp82_out1;
reg [7:0] cmp82_in0;
reg [7:0] cmp82_in1;

//-------dec layer:5----------
wire [7:0] cmp83_out0;
wire [7:0] cmp83_out1;
reg [7:0] cmp83_in0;
reg [7:0] cmp83_in1;

wire [7:0] cmp84_out0;
wire [7:0] cmp84_out1;
reg [7:0] cmp84_in0;
reg [7:0] cmp84_in1;

wire [7:0] cmp85_out0;
wire [7:0] cmp85_out1;
reg [7:0] cmp85_in0;
reg [7:0] cmp85_in1;

wire [7:0] cmp86_out0;
wire [7:0] cmp86_out1;
reg [7:0] cmp86_in0;
reg [7:0] cmp86_in1;

wire [7:0] cmp87_out0;
wire [7:0] cmp87_out1;
reg [7:0] cmp87_in0;
reg [7:0] cmp87_in1;

wire [7:0] cmp88_out0;
wire [7:0] cmp88_out1;
reg [7:0] cmp88_in0;
reg [7:0] cmp88_in1;

wire [7:0] cmp89_out0;
wire [7:0] cmp89_out1;
reg [7:0] cmp89_in0;
reg [7:0] cmp89_in1;

wire [7:0] cmp90_out0;
wire [7:0] cmp90_out1;
reg [7:0] cmp90_in0;
reg [7:0] cmp90_in1;

wire [7:0] cmp91_out0;
wire [7:0] cmp91_out1;
reg [7:0] cmp91_in0;
reg [7:0] cmp91_in1;

wire [7:0] cmp92_out0;
wire [7:0] cmp92_out1;
reg [7:0] cmp92_in0;
reg [7:0] cmp92_in1;

wire [7:0] cmp93_out0;
wire [7:0] cmp93_out1;
reg [7:0] cmp93_in0;
reg [7:0] cmp93_in1;

wire [7:0] cmp94_out0;
wire [7:0] cmp94_out1;
reg [7:0] cmp94_in0;
reg [7:0] cmp94_in1;

wire [7:0] cmp95_out0;
wire [7:0] cmp95_out1;
reg [7:0] cmp95_in0;
reg [7:0] cmp95_in1;

wire [7:0] cmp96_out0;
wire [7:0] cmp96_out1;
reg [7:0] cmp96_in0;
reg [7:0] cmp96_in1;

wire [7:0] cmp97_out0;
wire [7:0] cmp97_out1;
reg [7:0] cmp97_in0;
reg [7:0] cmp97_in1;

wire [7:0] cmp98_out0;
wire [7:0] cmp98_out1;
reg [7:0] cmp98_in0;
reg [7:0] cmp98_in1;

wire [7:0] cmp99_out0;
wire [7:0] cmp99_out1;
reg [7:0] cmp99_in0;
reg [7:0] cmp99_in1;

wire [7:0] cmp100_out0;
wire [7:0] cmp100_out1;
reg [7:0] cmp100_in0;
reg [7:0] cmp100_in1;

wire [7:0] cmp101_out0;
wire [7:0] cmp101_out1;
reg [7:0] cmp101_in0;
reg [7:0] cmp101_in1;

wire [7:0] cmp102_out0;
wire [7:0] cmp102_out1;
reg [7:0] cmp102_in0;
reg [7:0] cmp102_in1;

wire [7:0] cmp103_out0;
wire [7:0] cmp103_out1;
reg [7:0] cmp103_in0;
reg [7:0] cmp103_in1;

//-------dec layer:6----------
wire [7:0] cmp104_out0;
wire [7:0] cmp104_out1;
reg [7:0] cmp104_in0;
reg [7:0] cmp104_in1;

wire [7:0] cmp105_out0;
wire [7:0] cmp105_out1;
reg [7:0] cmp105_in0;
reg [7:0] cmp105_in1;

wire [7:0] cmp106_out0;
wire [7:0] cmp106_out1;
reg [7:0] cmp106_in0;
reg [7:0] cmp106_in1;

wire [7:0] cmp107_out0;
wire [7:0] cmp107_out1;
reg [7:0] cmp107_in0;
reg [7:0] cmp107_in1;

wire [7:0] cmp108_out0;
wire [7:0] cmp108_out1;
reg [7:0] cmp108_in0;
reg [7:0] cmp108_in1;

wire [7:0] cmp109_out0;
wire [7:0] cmp109_out1;
reg [7:0] cmp109_in0;
reg [7:0] cmp109_in1;

wire [7:0] cmp110_out0;
wire [7:0] cmp110_out1;
reg [7:0] cmp110_in0;
reg [7:0] cmp110_in1;

wire [7:0] cmp111_out0;
wire [7:0] cmp111_out1;
reg [7:0] cmp111_in0;
reg [7:0] cmp111_in1;

wire [7:0] cmp112_out0;
wire [7:0] cmp112_out1;
reg [7:0] cmp112_in0;
reg [7:0] cmp112_in1;

wire [7:0] cmp113_out0;
wire [7:0] cmp113_out1;
reg [7:0] cmp113_in0;
reg [7:0] cmp113_in1;

wire [7:0] cmp114_out0;
wire [7:0] cmp114_out1;
reg [7:0] cmp114_in0;
reg [7:0] cmp114_in1;

wire [7:0] cmp115_out0;
wire [7:0] cmp115_out1;
reg [7:0] cmp115_in0;
reg [7:0] cmp115_in1;

wire [7:0] cmp116_out0;
wire [7:0] cmp116_out1;
reg [7:0] cmp116_in0;
reg [7:0] cmp116_in1;

wire [7:0] cmp117_out0;
wire [7:0] cmp117_out1;
reg [7:0] cmp117_in0;
reg [7:0] cmp117_in1;

wire [7:0] cmp118_out0;
wire [7:0] cmp118_out1;
reg [7:0] cmp118_in0;
reg [7:0] cmp118_in1;

wire [7:0] cmp119_out0;
wire [7:0] cmp119_out1;
reg [7:0] cmp119_in0;
reg [7:0] cmp119_in1;

wire [7:0] cmp120_out0;
wire [7:0] cmp120_out1;
reg [7:0] cmp120_in0;
reg [7:0] cmp120_in1;

wire [7:0] cmp121_out0;
wire [7:0] cmp121_out1;
reg [7:0] cmp121_in0;
reg [7:0] cmp121_in1;

wire [7:0] cmp122_out0;
wire [7:0] cmp122_out1;
reg [7:0] cmp122_in0;
reg [7:0] cmp122_in1;

wire [7:0] cmp123_out0;
wire [7:0] cmp123_out1;
reg [7:0] cmp123_in0;
reg [7:0] cmp123_in1;

//-------dec layer:7----------
wire [7:0] cmp124_out0;
wire [7:0] cmp124_out1;
reg [7:0] cmp124_in0;
reg [7:0] cmp124_in1;

wire [7:0] cmp125_out0;
wire [7:0] cmp125_out1;
reg [7:0] cmp125_in0;
reg [7:0] cmp125_in1;

wire [7:0] cmp126_out0;
wire [7:0] cmp126_out1;
reg [7:0] cmp126_in0;
reg [7:0] cmp126_in1;

wire [7:0] cmp127_out0;
wire [7:0] cmp127_out1;
reg [7:0] cmp127_in0;
reg [7:0] cmp127_in1;

wire [7:0] cmp128_out0;
wire [7:0] cmp128_out1;
reg [7:0] cmp128_in0;
reg [7:0] cmp128_in1;

wire [7:0] cmp129_out0;
wire [7:0] cmp129_out1;
reg [7:0] cmp129_in0;
reg [7:0] cmp129_in1;

wire [7:0] cmp130_out0;
wire [7:0] cmp130_out1;
reg [7:0] cmp130_in0;
reg [7:0] cmp130_in1;

wire [7:0] cmp131_out0;
wire [7:0] cmp131_out1;
reg [7:0] cmp131_in0;
reg [7:0] cmp131_in1;

wire [7:0] cmp132_out0;
wire [7:0] cmp132_out1;
reg [7:0] cmp132_in0;
reg [7:0] cmp132_in1;

//-------dec layer:8----------
wire [7:0] cmp133_out0;
wire [7:0] cmp133_out1;
reg [7:0] cmp133_in0;
reg [7:0] cmp133_in1;

wire [7:0] cmp134_out0;
wire [7:0] cmp134_out1;
reg [7:0] cmp134_in0;
reg [7:0] cmp134_in1;

wire [7:0] cmp135_out0;
wire [7:0] cmp135_out1;
reg [7:0] cmp135_in0;
reg [7:0] cmp135_in1;

wire [7:0] cmp136_out0;
wire [7:0] cmp136_out1;
reg [7:0] cmp136_in0;
reg [7:0] cmp136_in1;

wire [7:0] cmp137_out0;
wire [7:0] cmp137_out1;
reg [7:0] cmp137_in0;
reg [7:0] cmp137_in1;

wire [7:0] cmp138_out0;
wire [7:0] cmp138_out1;
reg [7:0] cmp138_in0;
reg [7:0] cmp138_in1;

wire [7:0] cmp139_out0;
wire [7:0] cmp139_out1;
reg [7:0] cmp139_in0;
reg [7:0] cmp139_in1;

wire [7:0] cmp140_out0;
wire [7:0] cmp140_out1;
reg [7:0] cmp140_in0;
reg [7:0] cmp140_in1;

wire [7:0] cmp141_out0;
wire [7:0] cmp141_out1;
reg [7:0] cmp141_in0;
reg [7:0] cmp141_in1;

wire [7:0] cmp142_out0;
wire [7:0] cmp142_out1;
reg [7:0] cmp142_in0;
reg [7:0] cmp142_in1;

wire [7:0] cmp143_out0;
wire [7:0] cmp143_out1;
reg [7:0] cmp143_in0;
reg [7:0] cmp143_in1;

wire [7:0] cmp144_out0;
wire [7:0] cmp144_out1;
reg [7:0] cmp144_in0;
reg [7:0] cmp144_in1;

wire [7:0] cmp145_out0;
wire [7:0] cmp145_out1;
reg [7:0] cmp145_in0;
reg [7:0] cmp145_in1;

wire [7:0] cmp146_out0;
wire [7:0] cmp146_out1;
reg [7:0] cmp146_in0;
reg [7:0] cmp146_in1;

wire [7:0] cmp147_out0;
wire [7:0] cmp147_out1;
reg [7:0] cmp147_in0;
reg [7:0] cmp147_in1;

wire [7:0] cmp148_out0;
wire [7:0] cmp148_out1;
reg [7:0] cmp148_in0;
reg [7:0] cmp148_in1;

wire [7:0] cmp149_out0;
wire [7:0] cmp149_out1;
reg [7:0] cmp149_in0;
reg [7:0] cmp149_in1;

//-------dec layer:9----------
wire [7:0] cmp150_out0;
wire [7:0] cmp150_out1;
reg [7:0] cmp150_in0;
reg [7:0] cmp150_in1;

wire [7:0] cmp151_out0;
wire [7:0] cmp151_out1;
reg [7:0] cmp151_in0;
reg [7:0] cmp151_in1;

wire [7:0] cmp152_out0;
wire [7:0] cmp152_out1;
reg [7:0] cmp152_in0;
reg [7:0] cmp152_in1;

wire [7:0] cmp153_out0;
wire [7:0] cmp153_out1;
reg [7:0] cmp153_in0;
reg [7:0] cmp153_in1;

wire [7:0] cmp154_out0;
wire [7:0] cmp154_out1;
reg [7:0] cmp154_in0;
reg [7:0] cmp154_in1;

wire [7:0] cmp155_out0;
wire [7:0] cmp155_out1;
reg [7:0] cmp155_in0;
reg [7:0] cmp155_in1;

wire [7:0] cmp156_out0;
wire [7:0] cmp156_out1;
reg [7:0] cmp156_in0;
reg [7:0] cmp156_in1;

wire [7:0] cmp157_out0;
wire [7:0] cmp157_out1;
reg [7:0] cmp157_in0;
reg [7:0] cmp157_in1;

wire [7:0] cmp158_out0;
wire [7:0] cmp158_out1;
reg [7:0] cmp158_in0;
reg [7:0] cmp158_in1;

wire [7:0] cmp159_out0;
wire [7:0] cmp159_out1;
reg [7:0] cmp159_in0;
reg [7:0] cmp159_in1;

wire [7:0] cmp160_out0;
wire [7:0] cmp160_out1;
reg [7:0] cmp160_in0;
reg [7:0] cmp160_in1;

wire [7:0] cmp161_out0;
wire [7:0] cmp161_out1;
reg [7:0] cmp161_in0;
reg [7:0] cmp161_in1;

wire [7:0] cmp162_out0;
wire [7:0] cmp162_out1;
reg [7:0] cmp162_in0;
reg [7:0] cmp162_in1;

wire [7:0] cmp163_out0;
wire [7:0] cmp163_out1;
reg [7:0] cmp163_in0;
reg [7:0] cmp163_in1;

wire [7:0] cmp164_out0;
wire [7:0] cmp164_out1;
reg [7:0] cmp164_in0;
reg [7:0] cmp164_in1;

wire [7:0] cmp165_out0;
wire [7:0] cmp165_out1;
reg [7:0] cmp165_in0;
reg [7:0] cmp165_in1;

wire [7:0] cmp166_out0;
wire [7:0] cmp166_out1;
reg [7:0] cmp166_in0;
reg [7:0] cmp166_in1;

wire [7:0] cmp167_out0;
wire [7:0] cmp167_out1;
reg [7:0] cmp167_in0;
reg [7:0] cmp167_in1;

wire [7:0] cmp168_out0;
wire [7:0] cmp168_out1;
reg [7:0] cmp168_in0;
reg [7:0] cmp168_in1;

wire [7:0] cmp169_out0;
wire [7:0] cmp169_out1;
reg [7:0] cmp169_in0;
reg [7:0] cmp169_in1;

wire [7:0] cmp170_out0;
wire [7:0] cmp170_out1;
reg [7:0] cmp170_in0;
reg [7:0] cmp170_in1;

wire [7:0] cmp171_out0;
wire [7:0] cmp171_out1;
reg [7:0] cmp171_in0;
reg [7:0] cmp171_in1;

wire [7:0] cmp172_out0;
wire [7:0] cmp172_out1;
reg [7:0] cmp172_in0;
reg [7:0] cmp172_in1;

//-------dec layer:10----------
wire [7:0] cmp173_out0;
wire [7:0] cmp173_out1;
reg [7:0] cmp173_in0;
reg [7:0] cmp173_in1;

wire [7:0] cmp174_out0;
wire [7:0] cmp174_out1;
reg [7:0] cmp174_in0;
reg [7:0] cmp174_in1;

wire [7:0] cmp175_out0;
wire [7:0] cmp175_out1;
reg [7:0] cmp175_in0;
reg [7:0] cmp175_in1;

wire [7:0] cmp176_out0;
wire [7:0] cmp176_out1;
reg [7:0] cmp176_in0;
reg [7:0] cmp176_in1;

wire [7:0] cmp177_out0;
wire [7:0] cmp177_out1;
reg [7:0] cmp177_in0;
reg [7:0] cmp177_in1;

wire [7:0] cmp178_out0;
wire [7:0] cmp178_out1;
reg [7:0] cmp178_in0;
reg [7:0] cmp178_in1;

wire [7:0] cmp179_out0;
wire [7:0] cmp179_out1;
reg [7:0] cmp179_in0;
reg [7:0] cmp179_in1;

wire [7:0] cmp180_out0;
wire [7:0] cmp180_out1;
reg [7:0] cmp180_in0;
reg [7:0] cmp180_in1;

wire [7:0] cmp181_out0;
wire [7:0] cmp181_out1;
reg [7:0] cmp181_in0;
reg [7:0] cmp181_in1;

wire [7:0] cmp182_out0;
wire [7:0] cmp182_out1;
reg [7:0] cmp182_in0;
reg [7:0] cmp182_in1;

wire [7:0] cmp183_out0;
wire [7:0] cmp183_out1;
reg [7:0] cmp183_in0;
reg [7:0] cmp183_in1;

wire [7:0] cmp184_out0;
wire [7:0] cmp184_out1;
reg [7:0] cmp184_in0;
reg [7:0] cmp184_in1;

wire [7:0] cmp185_out0;
wire [7:0] cmp185_out1;
reg [7:0] cmp185_in0;
reg [7:0] cmp185_in1;

wire [7:0] cmp186_out0;
wire [7:0] cmp186_out1;
reg [7:0] cmp186_in0;
reg [7:0] cmp186_in1;

wire [7:0] cmp187_out0;
wire [7:0] cmp187_out1;
reg [7:0] cmp187_in0;
reg [7:0] cmp187_in1;

wire [7:0] cmp188_out0;
wire [7:0] cmp188_out1;
reg [7:0] cmp188_in0;
reg [7:0] cmp188_in1;

wire [7:0] cmp189_out0;
wire [7:0] cmp189_out1;
reg [7:0] cmp189_in0;
reg [7:0] cmp189_in1;

wire [7:0] cmp190_out0;
wire [7:0] cmp190_out1;
reg [7:0] cmp190_in0;
reg [7:0] cmp190_in1;

wire [7:0] cmp191_out0;
wire [7:0] cmp191_out1;
reg [7:0] cmp191_in0;
reg [7:0] cmp191_in1;

wire [7:0] cmp192_out0;
wire [7:0] cmp192_out1;
reg [7:0] cmp192_in0;
reg [7:0] cmp192_in1;

wire [7:0] cmp193_out0;
wire [7:0] cmp193_out1;
reg [7:0] cmp193_in0;
reg [7:0] cmp193_in1;

wire [7:0] cmp194_out0;
wire [7:0] cmp194_out1;
reg [7:0] cmp194_in0;
reg [7:0] cmp194_in1;

//-------dec layer:11----------
wire [7:0] cmp195_out0;
wire [7:0] cmp195_out1;
reg [7:0] cmp195_in0;
reg [7:0] cmp195_in1;

wire [7:0] cmp196_out0;
wire [7:0] cmp196_out1;
reg [7:0] cmp196_in0;
reg [7:0] cmp196_in1;

wire [7:0] cmp197_out0;
wire [7:0] cmp197_out1;
reg [7:0] cmp197_in0;
reg [7:0] cmp197_in1;

wire [7:0] cmp198_out0;
wire [7:0] cmp198_out1;
reg [7:0] cmp198_in0;
reg [7:0] cmp198_in1;

wire [7:0] cmp199_out0;
wire [7:0] cmp199_out1;
reg [7:0] cmp199_in0;
reg [7:0] cmp199_in1;

wire [7:0] cmp200_out0;
wire [7:0] cmp200_out1;
reg [7:0] cmp200_in0;
reg [7:0] cmp200_in1;

wire [7:0] cmp201_out0;
wire [7:0] cmp201_out1;
reg [7:0] cmp201_in0;
reg [7:0] cmp201_in1;

wire [7:0] cmp202_out0;
wire [7:0] cmp202_out1;
reg [7:0] cmp202_in0;
reg [7:0] cmp202_in1;

wire [7:0] cmp203_out0;
wire [7:0] cmp203_out1;
reg [7:0] cmp203_in0;
reg [7:0] cmp203_in1;

//-------dec layer:12----------
wire [7:0] cmp204_out0;
wire [7:0] cmp204_out1;
reg [7:0] cmp204_in0;
reg [7:0] cmp204_in1;

wire [7:0] cmp205_out0;
wire [7:0] cmp205_out1;
reg [7:0] cmp205_in0;
reg [7:0] cmp205_in1;

wire [7:0] cmp206_out0;
wire [7:0] cmp206_out1;
reg [7:0] cmp206_in0;
reg [7:0] cmp206_in1;

wire [7:0] cmp207_out0;
wire [7:0] cmp207_out1;
reg [7:0] cmp207_in0;
reg [7:0] cmp207_in1;

wire [7:0] cmp208_out0;
wire [7:0] cmp208_out1;
reg [7:0] cmp208_in0;
reg [7:0] cmp208_in1;

wire [7:0] cmp209_out0;
wire [7:0] cmp209_out1;
reg [7:0] cmp209_in0;
reg [7:0] cmp209_in1;

wire [7:0] cmp210_out0;
wire [7:0] cmp210_out1;
reg [7:0] cmp210_in0;
reg [7:0] cmp210_in1;

wire [7:0] cmp211_out0;
wire [7:0] cmp211_out1;
reg [7:0] cmp211_in0;
reg [7:0] cmp211_in1;

wire [7:0] cmp212_out0;
wire [7:0] cmp212_out1;
reg [7:0] cmp212_in0;
reg [7:0] cmp212_in1;

wire [7:0] cmp213_out0;
wire [7:0] cmp213_out1;
reg [7:0] cmp213_in0;
reg [7:0] cmp213_in1;

wire [7:0] cmp214_out0;
wire [7:0] cmp214_out1;
reg [7:0] cmp214_in0;
reg [7:0] cmp214_in1;

wire [7:0] cmp215_out0;
wire [7:0] cmp215_out1;
reg [7:0] cmp215_in0;
reg [7:0] cmp215_in1;

wire [7:0] cmp216_out0;
wire [7:0] cmp216_out1;
reg [7:0] cmp216_in0;
reg [7:0] cmp216_in1;

wire [7:0] cmp217_out0;
wire [7:0] cmp217_out1;
reg [7:0] cmp217_in0;
reg [7:0] cmp217_in1;

wire [7:0] cmp218_out0;
wire [7:0] cmp218_out1;
reg [7:0] cmp218_in0;
reg [7:0] cmp218_in1;

wire [7:0] cmp219_out0;
wire [7:0] cmp219_out1;
reg [7:0] cmp219_in0;
reg [7:0] cmp219_in1;

wire [7:0] cmp220_out0;
wire [7:0] cmp220_out1;
reg [7:0] cmp220_in0;
reg [7:0] cmp220_in1;

//-------dec layer:13----------
wire [7:0] cmp221_out0;
wire [7:0] cmp221_out1;
reg [7:0] cmp221_in0;
reg [7:0] cmp221_in1;

wire [7:0] cmp222_out0;
wire [7:0] cmp222_out1;
reg [7:0] cmp222_in0;
reg [7:0] cmp222_in1;

wire [7:0] cmp223_out0;
wire [7:0] cmp223_out1;
reg [7:0] cmp223_in0;
reg [7:0] cmp223_in1;

wire [7:0] cmp224_out0;
wire [7:0] cmp224_out1;
reg [7:0] cmp224_in0;
reg [7:0] cmp224_in1;

wire [7:0] cmp225_out0;
wire [7:0] cmp225_out1;
reg [7:0] cmp225_in0;
reg [7:0] cmp225_in1;

wire [7:0] cmp226_out0;
wire [7:0] cmp226_out1;
reg [7:0] cmp226_in0;
reg [7:0] cmp226_in1;

wire [7:0] cmp227_out0;
wire [7:0] cmp227_out1;
reg [7:0] cmp227_in0;
reg [7:0] cmp227_in1;

wire [7:0] cmp228_out0;
wire [7:0] cmp228_out1;
reg [7:0] cmp228_in0;
reg [7:0] cmp228_in1;

wire [7:0] cmp229_out0;
wire [7:0] cmp229_out1;
reg [7:0] cmp229_in0;
reg [7:0] cmp229_in1;

wire [7:0] cmp230_out0;
wire [7:0] cmp230_out1;
reg [7:0] cmp230_in0;
reg [7:0] cmp230_in1;

wire [7:0] cmp231_out0;
wire [7:0] cmp231_out1;
reg [7:0] cmp231_in0;
reg [7:0] cmp231_in1;

wire [7:0] cmp232_out0;
wire [7:0] cmp232_out1;
reg [7:0] cmp232_in0;
reg [7:0] cmp232_in1;

wire [7:0] cmp233_out0;
wire [7:0] cmp233_out1;
reg [7:0] cmp233_in0;
reg [7:0] cmp233_in1;

wire [7:0] cmp234_out0;
wire [7:0] cmp234_out1;
reg [7:0] cmp234_in0;
reg [7:0] cmp234_in1;

wire [7:0] cmp235_out0;
wire [7:0] cmp235_out1;
reg [7:0] cmp235_in0;
reg [7:0] cmp235_in1;

wire [7:0] cmp236_out0;
wire [7:0] cmp236_out1;
reg [7:0] cmp236_in0;
reg [7:0] cmp236_in1;

wire [7:0] cmp237_out0;
wire [7:0] cmp237_out1;
reg [7:0] cmp237_in0;
reg [7:0] cmp237_in1;

wire [7:0] cmp238_out0;
wire [7:0] cmp238_out1;
reg [7:0] cmp238_in0;
reg [7:0] cmp238_in1;

wire [7:0] cmp239_out0;
wire [7:0] cmp239_out1;
reg [7:0] cmp239_in0;
reg [7:0] cmp239_in1;

wire [7:0] cmp240_out0;
wire [7:0] cmp240_out1;
reg [7:0] cmp240_in0;
reg [7:0] cmp240_in1;

wire [7:0] cmp241_out0;
wire [7:0] cmp241_out1;
reg [7:0] cmp241_in0;
reg [7:0] cmp241_in1;

//-------dec layer:14----------
wire [7:0] cmp242_out0;
wire [7:0] cmp242_out1;
reg [7:0] cmp242_in0;
reg [7:0] cmp242_in1;

wire [7:0] cmp243_out0;
wire [7:0] cmp243_out1;
reg [7:0] cmp243_in0;
reg [7:0] cmp243_in1;

wire [7:0] cmp244_out0;
wire [7:0] cmp244_out1;
reg [7:0] cmp244_in0;
reg [7:0] cmp244_in1;

wire [7:0] cmp245_out0;
wire [7:0] cmp245_out1;
reg [7:0] cmp245_in0;
reg [7:0] cmp245_in1;

wire [7:0] cmp246_out0;
wire [7:0] cmp246_out1;
reg [7:0] cmp246_in0;
reg [7:0] cmp246_in1;

wire [7:0] cmp247_out0;
wire [7:0] cmp247_out1;
reg [7:0] cmp247_in0;
reg [7:0] cmp247_in1;

wire [7:0] cmp248_out0;
wire [7:0] cmp248_out1;
reg [7:0] cmp248_in0;
reg [7:0] cmp248_in1;

wire [7:0] cmp249_out0;
wire [7:0] cmp249_out1;
reg [7:0] cmp249_in0;
reg [7:0] cmp249_in1;

wire [7:0] cmp250_out0;
wire [7:0] cmp250_out1;
reg [7:0] cmp250_in0;
reg [7:0] cmp250_in1;

wire [7:0] cmp251_out0;
wire [7:0] cmp251_out1;
reg [7:0] cmp251_in0;
reg [7:0] cmp251_in1;

wire [7:0] cmp252_out0;
wire [7:0] cmp252_out1;
reg [7:0] cmp252_in0;
reg [7:0] cmp252_in1;

wire [7:0] cmp253_out0;
wire [7:0] cmp253_out1;
reg [7:0] cmp253_in0;
reg [7:0] cmp253_in1;

wire [7:0] cmp254_out0;
wire [7:0] cmp254_out1;
reg [7:0] cmp254_in0;
reg [7:0] cmp254_in1;

wire [7:0] cmp255_out0;
wire [7:0] cmp255_out1;
reg [7:0] cmp255_in0;
reg [7:0] cmp255_in1;

wire [7:0] cmp256_out0;
wire [7:0] cmp256_out1;
reg [7:0] cmp256_in0;
reg [7:0] cmp256_in1;

wire [7:0] cmp257_out0;
wire [7:0] cmp257_out1;
reg [7:0] cmp257_in0;
reg [7:0] cmp257_in1;

wire [7:0] cmp258_out0;
wire [7:0] cmp258_out1;
reg [7:0] cmp258_in0;
reg [7:0] cmp258_in1;

wire [7:0] cmp259_out0;
wire [7:0] cmp259_out1;
reg [7:0] cmp259_in0;
reg [7:0] cmp259_in1;

wire [7:0] cmp260_out0;
wire [7:0] cmp260_out1;
reg [7:0] cmp260_in0;
reg [7:0] cmp260_in1;

wire [7:0] cmp261_out0;
wire [7:0] cmp261_out1;
reg [7:0] cmp261_in0;
reg [7:0] cmp261_in1;

wire [7:0] cmp262_out0;
wire [7:0] cmp262_out1;
reg [7:0] cmp262_in0;
reg [7:0] cmp262_in1;

wire [7:0] cmp263_out0;
wire [7:0] cmp263_out1;
reg [7:0] cmp263_in0;
reg [7:0] cmp263_in1;

wire [7:0] cmp264_out0;
wire [7:0] cmp264_out1;
reg [7:0] cmp264_in0;
reg [7:0] cmp264_in1;

wire [7:0] cmp265_out0;
wire [7:0] cmp265_out1;
reg [7:0] cmp265_in0;
reg [7:0] cmp265_in1;

//-------dec layer:15----------
wire [7:0] cmp266_out0;
wire [7:0] cmp266_out1;
reg [7:0] cmp266_in0;
reg [7:0] cmp266_in1;

wire [7:0] cmp267_out0;
wire [7:0] cmp267_out1;
reg [7:0] cmp267_in0;
reg [7:0] cmp267_in1;

wire [7:0] cmp268_out0;
wire [7:0] cmp268_out1;
reg [7:0] cmp268_in0;
reg [7:0] cmp268_in1;

wire [7:0] cmp269_out0;
wire [7:0] cmp269_out1;
reg [7:0] cmp269_in0;
reg [7:0] cmp269_in1;

wire [7:0] cmp270_out0;
wire [7:0] cmp270_out1;
reg [7:0] cmp270_in0;
reg [7:0] cmp270_in1;

wire [7:0] cmp271_out0;
wire [7:0] cmp271_out1;
reg [7:0] cmp271_in0;
reg [7:0] cmp271_in1;

wire [7:0] cmp272_out0;
wire [7:0] cmp272_out1;
reg [7:0] cmp272_in0;
reg [7:0] cmp272_in1;

wire [7:0] cmp273_out0;
wire [7:0] cmp273_out1;
reg [7:0] cmp273_in0;
reg [7:0] cmp273_in1;

wire [7:0] cmp274_out0;
wire [7:0] cmp274_out1;
reg [7:0] cmp274_in0;
reg [7:0] cmp274_in1;

wire [7:0] cmp275_out0;
wire [7:0] cmp275_out1;
reg [7:0] cmp275_in0;
reg [7:0] cmp275_in1;

wire [7:0] cmp276_out0;
wire [7:0] cmp276_out1;
reg [7:0] cmp276_in0;
reg [7:0] cmp276_in1;

wire [7:0] cmp277_out0;
wire [7:0] cmp277_out1;
reg [7:0] cmp277_in0;
reg [7:0] cmp277_in1;

wire [7:0] cmp278_out0;
wire [7:0] cmp278_out1;
reg [7:0] cmp278_in0;
reg [7:0] cmp278_in1;

wire [7:0] cmp279_out0;
wire [7:0] cmp279_out1;
reg [7:0] cmp279_in0;
reg [7:0] cmp279_in1;

wire [7:0] cmp280_out0;
wire [7:0] cmp280_out1;
reg [7:0] cmp280_in0;
reg [7:0] cmp280_in1;

wire [7:0] cmp281_out0;
wire [7:0] cmp281_out1;
reg [7:0] cmp281_in0;
reg [7:0] cmp281_in1;

wire [7:0] cmp282_out0;
wire [7:0] cmp282_out1;
reg [7:0] cmp282_in0;
reg [7:0] cmp282_in1;

wire [7:0] cmp283_out0;
wire [7:0] cmp283_out1;
reg [7:0] cmp283_in0;
reg [7:0] cmp283_in1;

wire [7:0] cmp284_out0;
wire [7:0] cmp284_out1;
reg [7:0] cmp284_in0;
reg [7:0] cmp284_in1;

wire [7:0] cmp285_out0;
wire [7:0] cmp285_out1;
reg [7:0] cmp285_in0;
reg [7:0] cmp285_in1;

wire [7:0] cmp286_out0;
wire [7:0] cmp286_out1;
reg [7:0] cmp286_in0;
reg [7:0] cmp286_in1;

wire [7:0] cmp287_out0;
wire [7:0] cmp287_out1;
reg [7:0] cmp287_in0;
reg [7:0] cmp287_in1;

wire [7:0] cmp288_out0;
wire [7:0] cmp288_out1;
reg [7:0] cmp288_in0;
reg [7:0] cmp288_in1;

//-------dec layer:16----------
wire [7:0] cmp289_out0;
wire [7:0] cmp289_out1;
reg [7:0] cmp289_in0;
reg [7:0] cmp289_in1;

wire [7:0] cmp290_out0;
wire [7:0] cmp290_out1;
reg [7:0] cmp290_in0;
reg [7:0] cmp290_in1;

wire [7:0] cmp291_out0;
wire [7:0] cmp291_out1;
reg [7:0] cmp291_in0;
reg [7:0] cmp291_in1;

wire [7:0] cmp292_out0;
wire [7:0] cmp292_out1;
reg [7:0] cmp292_in0;
reg [7:0] cmp292_in1;

wire [7:0] cmp293_out0;
wire [7:0] cmp293_out1;
reg [7:0] cmp293_in0;
reg [7:0] cmp293_in1;

wire [7:0] cmp294_out0;
wire [7:0] cmp294_out1;
reg [7:0] cmp294_in0;
reg [7:0] cmp294_in1;

wire [7:0] cmp295_out0;
wire [7:0] cmp295_out1;
reg [7:0] cmp295_in0;
reg [7:0] cmp295_in1;

wire [7:0] cmp296_out0;
wire [7:0] cmp296_out1;
reg [7:0] cmp296_in0;
reg [7:0] cmp296_in1;

wire [7:0] cmp297_out0;
wire [7:0] cmp297_out1;
reg [7:0] cmp297_in0;
reg [7:0] cmp297_in1;

//-------dec layer:17----------
wire [7:0] cmp298_out0;
wire [7:0] cmp298_out1;
reg [7:0] cmp298_in0;
reg [7:0] cmp298_in1;

wire [7:0] cmp299_out0;
wire [7:0] cmp299_out1;
reg [7:0] cmp299_in0;
reg [7:0] cmp299_in1;

wire [7:0] cmp300_out0;
wire [7:0] cmp300_out1;
reg [7:0] cmp300_in0;
reg [7:0] cmp300_in1;

wire [7:0] cmp301_out0;
wire [7:0] cmp301_out1;
reg [7:0] cmp301_in0;
reg [7:0] cmp301_in1;

wire [7:0] cmp302_out0;
wire [7:0] cmp302_out1;
reg [7:0] cmp302_in0;
reg [7:0] cmp302_in1;

wire [7:0] cmp303_out0;
wire [7:0] cmp303_out1;
reg [7:0] cmp303_in0;
reg [7:0] cmp303_in1;

wire [7:0] cmp304_out0;
wire [7:0] cmp304_out1;
reg [7:0] cmp304_in0;
reg [7:0] cmp304_in1;

wire [7:0] cmp305_out0;
wire [7:0] cmp305_out1;
reg [7:0] cmp305_in0;
reg [7:0] cmp305_in1;

//-------dec layer:18----------
wire [7:0] cmp306_out0;
wire [7:0] cmp306_out1;
reg [7:0] cmp306_in0;
reg [7:0] cmp306_in1;

wire [7:0] cmp307_out0;
wire [7:0] cmp307_out1;
reg [7:0] cmp307_in0;
reg [7:0] cmp307_in1;

wire [7:0] cmp308_out0;
wire [7:0] cmp308_out1;
reg [7:0] cmp308_in0;
reg [7:0] cmp308_in1;

wire [7:0] cmp309_out0;
wire [7:0] cmp309_out1;
reg [7:0] cmp309_in0;
reg [7:0] cmp309_in1;

//-------dec layer:19----------
wire [7:0] cmp310_out0;
wire [7:0] cmp310_out1;
reg [7:0] cmp310_in0;
reg [7:0] cmp310_in1;

wire [7:0] cmp311_out0;
wire [7:0] cmp311_out1;
reg [7:0] cmp311_in0;
reg [7:0] cmp311_in1;

//-------dec layer:20----------
wire [7:0] cmp312_out0;
wire [7:0] cmp312_out1;
reg [7:0] cmp312_in0;
reg [7:0] cmp312_in1;

//-------Temp Register----------
reg [7:0] r_0_17_tmp;
reg [7:0] r_0_18_tmp;
reg [7:0] r_0_19_tmp;
reg [7:0] r_0_20_tmp;
reg [7:0] r_0_21_tmp;
reg [7:0] r_0_22_tmp;
reg [7:0] r_0_23_tmp;
reg [7:0] r_0_24_tmp;
reg [7:0] r_0_25_tmp;
reg [7:0] r_0_26_tmp;
reg [7:0] r_0_27_tmp;
reg [7:0] r_0_28_tmp;
reg [7:0] r_0_29_tmp;
reg [7:0] r_0_30_tmp;
reg [7:0] r_0_31_tmp;
reg [7:0] r_1_33_tmp;
reg [7:0] r_1_34_tmp;
reg [7:0] r_1_35_tmp;
reg [7:0] r_1_36_tmp;
reg [7:0] r_1_37_tmp;
reg [7:0] r_1_38_tmp;
reg [7:0] r_1_39_tmp;
reg [7:0] r_1_40_tmp;
reg [7:0] r_1_41_tmp;
reg [7:0] r_1_42_tmp;
reg [7:0] r_1_43_tmp;
reg [7:0] r_1_44_tmp;
reg [7:0] r_1_45_tmp;
reg [7:0] r_1_46_tmp;
reg [7:0] r_1_47_tmp;
reg [7:0] r_2_48_tmp;
reg [7:0] r_3_0_tmp;
reg [7:0] r_3_1_tmp;
reg [7:0] r_3_2_tmp;
reg [7:0] r_3_3_tmp;
reg [7:0] r_3_4_tmp;
reg [7:0] r_3_5_tmp;
reg [7:0] r_3_6_tmp;
reg [7:0] r_3_7_tmp;
reg [7:0] r_3_8_tmp;
reg [7:0] r_3_9_tmp;
reg [7:0] r_3_10_tmp;
reg [7:0] r_3_11_tmp;
reg [7:0] r_3_12_tmp;
reg [7:0] r_3_13_tmp;
reg [7:0] r_3_14_tmp;
reg [7:0] r_3_15_tmp;
reg [7:0] r_3_48_tmp;
reg [7:0] r_4_0_tmp;
reg [7:0] r_4_1_tmp;
reg [7:0] r_4_2_tmp;
reg [7:0] r_4_3_tmp;
reg [7:0] r_4_4_tmp;
reg [7:0] r_4_5_tmp;
reg [7:0] r_4_6_tmp;
reg [7:0] r_4_7_tmp;
reg [7:0] r_4_16_tmp;
reg [7:0] r_4_17_tmp;
reg [7:0] r_4_18_tmp;
reg [7:0] r_4_19_tmp;
reg [7:0] r_4_20_tmp;
reg [7:0] r_4_21_tmp;
reg [7:0] r_4_22_tmp;
reg [7:0] r_4_23_tmp;
reg [7:0] r_4_25_tmp;
reg [7:0] r_4_26_tmp;
reg [7:0] r_4_27_tmp;
reg [7:0] r_4_28_tmp;
reg [7:0] r_4_29_tmp;
reg [7:0] r_4_30_tmp;
reg [7:0] r_4_31_tmp;
reg [7:0] r_4_40_tmp;
reg [7:0] r_4_41_tmp;
reg [7:0] r_4_42_tmp;
reg [7:0] r_4_43_tmp;
reg [7:0] r_4_44_tmp;
reg [7:0] r_4_45_tmp;
reg [7:0] r_4_46_tmp;
reg [7:0] r_4_47_tmp;
reg [7:0] r_5_41_tmp;
reg [7:0] r_5_42_tmp;
reg [7:0] r_5_43_tmp;
reg [7:0] r_5_44_tmp;
reg [7:0] r_5_45_tmp;
reg [7:0] r_5_46_tmp;
reg [7:0] r_5_47_tmp;
reg [7:0] r_6_0_tmp;
reg [7:0] r_6_1_tmp;
reg [7:0] r_6_2_tmp;
reg [7:0] r_6_3_tmp;
reg [7:0] r_6_4_tmp;
reg [7:0] r_6_5_tmp;
reg [7:0] r_6_6_tmp;
reg [7:0] r_6_7_tmp;
reg [7:0] r_6_48_tmp;
reg [7:0] r_7_0_tmp;
reg [7:0] r_7_1_tmp;
reg [7:0] r_7_2_tmp;
reg [7:0] r_7_3_tmp;
reg [7:0] r_7_8_tmp;
reg [7:0] r_7_9_tmp;
reg [7:0] r_7_10_tmp;
reg [7:0] r_7_11_tmp;
reg [7:0] r_7_16_tmp;
reg [7:0] r_7_17_tmp;
reg [7:0] r_7_18_tmp;
reg [7:0] r_7_19_tmp;
reg [7:0] r_7_21_tmp;
reg [7:0] r_7_22_tmp;
reg [7:0] r_7_23_tmp;
reg [7:0] r_7_24_tmp;
reg [7:0] r_7_25_tmp;
reg [7:0] r_7_26_tmp;
reg [7:0] r_7_27_tmp;
reg [7:0] r_7_28_tmp;
reg [7:0] r_7_29_tmp;
reg [7:0] r_7_30_tmp;
reg [7:0] r_7_31_tmp;
reg [7:0] r_7_36_tmp;
reg [7:0] r_7_37_tmp;
reg [7:0] r_7_38_tmp;
reg [7:0] r_7_39_tmp;
reg [7:0] r_7_44_tmp;
reg [7:0] r_7_45_tmp;
reg [7:0] r_7_46_tmp;
reg [7:0] r_7_47_tmp;
reg [7:0] r_8_0_tmp;
reg [7:0] r_8_1_tmp;
reg [7:0] r_8_2_tmp;
reg [7:0] r_8_3_tmp;
reg [7:0] r_8_8_tmp;
reg [7:0] r_8_9_tmp;
reg [7:0] r_8_10_tmp;
reg [7:0] r_8_11_tmp;
reg [7:0] r_8_37_tmp;
reg [7:0] r_8_38_tmp;
reg [7:0] r_8_39_tmp;
reg [7:0] r_8_44_tmp;
reg [7:0] r_8_45_tmp;
reg [7:0] r_8_46_tmp;
reg [7:0] r_8_47_tmp;
reg [7:0] r_9_45_tmp;
reg [7:0] r_9_46_tmp;
reg [7:0] r_9_47_tmp;
reg [7:0] r_10_0_tmp;
reg [7:0] r_10_1_tmp;
reg [7:0] r_10_2_tmp;
reg [7:0] r_10_3_tmp;
reg [7:0] r_10_48_tmp;
reg [7:0] r_11_0_tmp;
reg [7:0] r_11_1_tmp;
reg [7:0] r_11_4_tmp;
reg [7:0] r_11_5_tmp;
reg [7:0] r_11_8_tmp;
reg [7:0] r_11_9_tmp;
reg [7:0] r_11_12_tmp;
reg [7:0] r_11_13_tmp;
reg [7:0] r_11_16_tmp;
reg [7:0] r_11_17_tmp;
reg [7:0] r_11_19_tmp;
reg [7:0] r_11_20_tmp;
reg [7:0] r_11_21_tmp;
reg [7:0] r_11_22_tmp;
reg [7:0] r_11_23_tmp;
reg [7:0] r_11_24_tmp;
reg [7:0] r_11_25_tmp;
reg [7:0] r_11_26_tmp;
reg [7:0] r_11_27_tmp;
reg [7:0] r_11_28_tmp;
reg [7:0] r_11_29_tmp;
reg [7:0] r_11_30_tmp;
reg [7:0] r_11_31_tmp;
reg [7:0] r_11_34_tmp;
reg [7:0] r_11_35_tmp;
reg [7:0] r_11_38_tmp;
reg [7:0] r_11_39_tmp;
reg [7:0] r_11_42_tmp;
reg [7:0] r_11_43_tmp;
reg [7:0] r_11_46_tmp;
reg [7:0] r_11_47_tmp;
reg [7:0] r_12_0_tmp;
reg [7:0] r_12_1_tmp;
reg [7:0] r_12_4_tmp;
reg [7:0] r_12_5_tmp;
reg [7:0] r_12_8_tmp;
reg [7:0] r_12_9_tmp;
reg [7:0] r_12_12_tmp;
reg [7:0] r_12_13_tmp;
reg [7:0] r_12_35_tmp;
reg [7:0] r_12_38_tmp;
reg [7:0] r_12_39_tmp;
reg [7:0] r_12_42_tmp;
reg [7:0] r_12_43_tmp;
reg [7:0] r_12_46_tmp;
reg [7:0] r_12_47_tmp;
reg [7:0] r_13_0_tmp;
reg [7:0] r_13_1_tmp;
reg [7:0] r_13_4_tmp;
reg [7:0] r_13_5_tmp;
reg [7:0] r_13_43_tmp;
reg [7:0] r_13_46_tmp;
reg [7:0] r_13_47_tmp;
reg [7:0] r_14_47_tmp;
reg [7:0] r_15_0_tmp;
reg [7:0] r_15_1_tmp;
reg [7:0] r_15_48_tmp;
reg [7:0] r_16_0_tmp;
reg [7:0] r_16_2_tmp;
reg [7:0] r_16_4_tmp;
reg [7:0] r_16_6_tmp;
reg [7:0] r_16_8_tmp;
reg [7:0] r_16_10_tmp;
reg [7:0] r_16_12_tmp;
reg [7:0] r_16_14_tmp;
reg [7:0] r_16_16_tmp;
reg [7:0] r_16_18_tmp;
reg [7:0] r_16_19_tmp;
reg [7:0] r_16_20_tmp;
reg [7:0] r_16_21_tmp;
reg [7:0] r_16_22_tmp;
reg [7:0] r_16_23_tmp;
reg [7:0] r_16_24_tmp;
reg [7:0] r_16_25_tmp;
reg [7:0] r_16_26_tmp;
reg [7:0] r_16_27_tmp;
reg [7:0] r_16_28_tmp;
reg [7:0] r_16_29_tmp;
reg [7:0] r_16_30_tmp;
reg [7:0] r_16_31_tmp;
reg [7:0] r_16_33_tmp;
reg [7:0] r_16_35_tmp;
reg [7:0] r_16_37_tmp;
reg [7:0] r_16_39_tmp;
reg [7:0] r_16_41_tmp;
reg [7:0] r_16_43_tmp;
reg [7:0] r_16_45_tmp;
reg [7:0] r_16_47_tmp;
reg [7:0] r_17_0_tmp;
reg [7:0] r_17_1_tmp;
reg [7:0] r_17_2_tmp;
reg [7:0] r_17_3_tmp;
reg [7:0] r_17_4_tmp;
reg [7:0] r_17_5_tmp;
reg [7:0] r_17_6_tmp;
reg [7:0] r_17_7_tmp;
reg [7:0] r_17_8_tmp;
reg [7:0] r_17_10_tmp;
reg [7:0] r_17_12_tmp;
reg [7:0] r_17_14_tmp;
reg [7:0] r_17_16_tmp;
reg [7:0] r_17_18_tmp;
reg [7:0] r_17_20_tmp;
reg [7:0] r_17_22_tmp;
reg [7:0] r_17_25_tmp;
reg [7:0] r_17_27_tmp;
reg [7:0] r_17_29_tmp;
reg [7:0] r_17_31_tmp;
reg [7:0] r_17_33_tmp;
reg [7:0] r_17_35_tmp;
reg [7:0] r_17_37_tmp;
reg [7:0] r_17_39_tmp;
reg [7:0] r_17_40_tmp;
reg [7:0] r_17_41_tmp;
reg [7:0] r_17_42_tmp;
reg [7:0] r_17_43_tmp;
reg [7:0] r_17_44_tmp;
reg [7:0] r_17_45_tmp;
reg [7:0] r_17_46_tmp;
reg [7:0] r_17_47_tmp;
reg [7:0] r_17_48_tmp;
reg [7:0] r_18_0_tmp;
reg [7:0] r_18_1_tmp;
reg [7:0] r_18_2_tmp;
reg [7:0] r_18_3_tmp;
reg [7:0] r_18_4_tmp;
reg [7:0] r_18_5_tmp;
reg [7:0] r_18_6_tmp;
reg [7:0] r_18_7_tmp;
reg [7:0] r_18_8_tmp;
reg [7:0] r_18_9_tmp;
reg [7:0] r_18_10_tmp;
reg [7:0] r_18_11_tmp;
reg [7:0] r_18_12_tmp;
reg [7:0] r_18_13_tmp;
reg [7:0] r_18_14_tmp;
reg [7:0] r_18_15_tmp;
reg [7:0] r_18_16_tmp;
reg [7:0] r_18_18_tmp;
reg [7:0] r_18_20_tmp;
reg [7:0] r_18_22_tmp;
reg [7:0] r_18_25_tmp;
reg [7:0] r_18_27_tmp;
reg [7:0] r_18_29_tmp;
reg [7:0] r_18_31_tmp;
reg [7:0] r_18_32_tmp;
reg [7:0] r_18_33_tmp;
reg [7:0] r_18_34_tmp;
reg [7:0] r_18_35_tmp;
reg [7:0] r_18_36_tmp;
reg [7:0] r_18_37_tmp;
reg [7:0] r_18_38_tmp;
reg [7:0] r_18_39_tmp;
reg [7:0] r_18_40_tmp;
reg [7:0] r_18_41_tmp;
reg [7:0] r_18_42_tmp;
reg [7:0] r_18_43_tmp;
reg [7:0] r_18_44_tmp;
reg [7:0] r_18_45_tmp;
reg [7:0] r_18_46_tmp;
reg [7:0] r_18_47_tmp;
reg [7:0] r_18_48_tmp;
reg [7:0] r_19_0_tmp;
reg [7:0] r_19_1_tmp;
reg [7:0] r_19_2_tmp;
reg [7:0] r_19_3_tmp;
reg [7:0] r_19_4_tmp;
reg [7:0] r_19_5_tmp;
reg [7:0] r_19_6_tmp;
reg [7:0] r_19_7_tmp;
reg [7:0] r_19_8_tmp;
reg [7:0] r_19_9_tmp;
reg [7:0] r_19_10_tmp;
reg [7:0] r_19_11_tmp;
reg [7:0] r_19_12_tmp;
reg [7:0] r_19_13_tmp;
reg [7:0] r_19_14_tmp;
reg [7:0] r_19_15_tmp;
reg [7:0] r_19_16_tmp;
reg [7:0] r_19_17_tmp;
reg [7:0] r_19_18_tmp;
reg [7:0] r_19_19_tmp;
reg [7:0] r_19_20_tmp;
reg [7:0] r_19_22_tmp;
reg [7:0] r_19_25_tmp;
reg [7:0] r_19_27_tmp;
reg [7:0] r_19_28_tmp;
reg [7:0] r_19_29_tmp;
reg [7:0] r_19_30_tmp;
reg [7:0] r_19_31_tmp;
reg [7:0] r_19_32_tmp;
reg [7:0] r_19_33_tmp;
reg [7:0] r_19_34_tmp;
reg [7:0] r_19_35_tmp;
reg [7:0] r_19_36_tmp;
reg [7:0] r_19_37_tmp;
reg [7:0] r_19_38_tmp;
reg [7:0] r_19_39_tmp;
reg [7:0] r_19_40_tmp;
reg [7:0] r_19_41_tmp;
reg [7:0] r_19_42_tmp;
reg [7:0] r_19_43_tmp;
reg [7:0] r_19_44_tmp;
reg [7:0] r_19_45_tmp;
reg [7:0] r_19_46_tmp;
reg [7:0] r_19_47_tmp;
reg [7:0] r_19_48_tmp;
reg [7:0] r_20_0_tmp;
reg [7:0] r_20_1_tmp;
reg [7:0] r_20_2_tmp;
reg [7:0] r_20_3_tmp;
reg [7:0] r_20_4_tmp;
reg [7:0] r_20_5_tmp;
reg [7:0] r_20_6_tmp;
reg [7:0] r_20_7_tmp;
reg [7:0] r_20_8_tmp;
reg [7:0] r_20_9_tmp;
reg [7:0] r_20_10_tmp;
reg [7:0] r_20_11_tmp;
reg [7:0] r_20_12_tmp;
reg [7:0] r_20_13_tmp;
reg [7:0] r_20_14_tmp;
reg [7:0] r_20_15_tmp;
reg [7:0] r_20_16_tmp;
reg [7:0] r_20_17_tmp;
reg [7:0] r_20_18_tmp;
reg [7:0] r_20_19_tmp;
reg [7:0] r_20_20_tmp;
reg [7:0] r_20_21_tmp;
reg [7:0] r_20_22_tmp;
reg [7:0] r_20_25_tmp;
reg [7:0] r_20_26_tmp;
reg [7:0] r_20_27_tmp;
reg [7:0] r_20_28_tmp;
reg [7:0] r_20_29_tmp;
reg [7:0] r_20_30_tmp;
reg [7:0] r_20_31_tmp;
reg [7:0] r_20_32_tmp;
reg [7:0] r_20_33_tmp;
reg [7:0] r_20_34_tmp;
reg [7:0] r_20_35_tmp;
reg [7:0] r_20_36_tmp;
reg [7:0] r_20_37_tmp;
reg [7:0] r_20_38_tmp;
reg [7:0] r_20_39_tmp;
reg [7:0] r_20_40_tmp;
reg [7:0] r_20_41_tmp;
reg [7:0] r_20_42_tmp;
reg [7:0] r_20_43_tmp;
reg [7:0] r_20_44_tmp;
reg [7:0] r_20_45_tmp;
reg [7:0] r_20_46_tmp;
reg [7:0] r_20_47_tmp;
reg [7:0] r_20_48_tmp;
//-----------------------------

always @(posedge clk)begin
//--------INPUT LAYER-------------
cmp0_in0 <= x_0;
cmp0_in1 <= x_32;
r0[0] <= cmp0_out0;
r0[32] <= cmp0_out1;

cmp1_in0 <= x_1;
cmp1_in1 <= x_33;
r0[1] <= cmp1_out0;
r0[33] <= cmp1_out1;

cmp2_in0 <= x_2;
cmp2_in1 <= x_34;
r0[2] <= cmp2_out0;
r0[34] <= cmp2_out1;

cmp3_in0 <= x_3;
cmp3_in1 <= x_35;
r0[3] <= cmp3_out0;
r0[35] <= cmp3_out1;

cmp4_in0 <= x_4;
cmp4_in1 <= x_36;
r0[4] <= cmp4_out0;
r0[36] <= cmp4_out1;

cmp5_in0 <= x_5;
cmp5_in1 <= x_37;
r0[5] <= cmp5_out0;
r0[37] <= cmp5_out1;

cmp6_in0 <= x_6;
cmp6_in1 <= x_38;
r0[6] <= cmp6_out0;
r0[38] <= cmp6_out1;

cmp7_in0 <= x_7;
cmp7_in1 <= x_39;
r0[7] <= cmp7_out0;
r0[39] <= cmp7_out1;

cmp8_in0 <= x_8;
cmp8_in1 <= x_40;
r0[8] <= cmp8_out0;
r0[40] <= cmp8_out1;

cmp9_in0 <= x_9;
cmp9_in1 <= x_41;
r0[9] <= cmp9_out0;
r0[41] <= cmp9_out1;

cmp10_in0 <= x_10;
cmp10_in1 <= x_42;
r0[10] <= cmp10_out0;
r0[42] <= cmp10_out1;

cmp11_in0 <= x_11;
cmp11_in1 <= x_43;
r0[11] <= cmp11_out0;
r0[43] <= cmp11_out1;

cmp12_in0 <= x_12;
cmp12_in1 <= x_44;
r0[12] <= cmp12_out0;
r0[44] <= cmp12_out1;

cmp13_in0 <= x_13;
cmp13_in1 <= x_45;
r0[13] <= cmp13_out0;
r0[45] <= cmp13_out1;

cmp14_in0 <= x_14;
cmp14_in1 <= x_46;
r0[14] <= cmp14_out0;
r0[46] <= cmp14_out1;

cmp15_in0 <= x_15;
cmp15_in1 <= x_47;
r0[15] <= cmp15_out0;
r0[47] <= cmp15_out1;

cmp16_in0 <= x_16;
cmp16_in1 <= x_48;
r0[16] <= cmp16_out0;
r0[48] <= cmp16_out1;

r_0_17_tmp <= x_17;
r0[17] <= r_0_17_tmp ;
r_0_18_tmp <= x_18;
r0[18] <= r_0_18_tmp ;
r_0_19_tmp <= x_19;
r0[19] <= r_0_19_tmp ;
r_0_20_tmp <= x_20;
r0[20] <= r_0_20_tmp ;
r_0_21_tmp <= x_21;
r0[21] <= r_0_21_tmp ;
r_0_22_tmp <= x_22;
r0[22] <= r_0_22_tmp ;
r_0_23_tmp <= x_23;
r0[23] <= r_0_23_tmp ;
r_0_24_tmp <= x_24;
r0[24] <= r_0_24_tmp ;
r_0_25_tmp <= x_25;
r0[25] <= r_0_25_tmp ;
r_0_26_tmp <= x_26;
r0[26] <= r_0_26_tmp ;
r_0_27_tmp <= x_27;
r0[27] <= r_0_27_tmp ;
r_0_28_tmp <= x_28;
r0[28] <= r_0_28_tmp ;
r_0_29_tmp <= x_29;
r0[29] <= r_0_29_tmp ;
r_0_30_tmp <= x_30;
r0[30] <= r_0_30_tmp ;
r_0_31_tmp <= x_31;
r0[31] <= r_0_31_tmp ;
//--------------------------

//---------layer : 1------------
cmp17_in0 <= r0[0];
cmp17_in1 <= r0[16];
r1[0] <= cmp17_out0;
r1[16] <= cmp17_out1;

cmp18_in0 <= r0[1];
cmp18_in1 <= r0[17];
r1[1] <= cmp18_out0;
r1[17] <= cmp18_out1;

cmp19_in0 <= r0[2];
cmp19_in1 <= r0[18];
r1[2] <= cmp19_out0;
r1[18] <= cmp19_out1;

cmp20_in0 <= r0[3];
cmp20_in1 <= r0[19];
r1[3] <= cmp20_out0;
r1[19] <= cmp20_out1;

cmp21_in0 <= r0[4];
cmp21_in1 <= r0[20];
r1[4] <= cmp21_out0;
r1[20] <= cmp21_out1;

cmp22_in0 <= r0[5];
cmp22_in1 <= r0[21];
r1[5] <= cmp22_out0;
r1[21] <= cmp22_out1;

cmp23_in0 <= r0[6];
cmp23_in1 <= r0[22];
r1[6] <= cmp23_out0;
r1[22] <= cmp23_out1;

cmp24_in0 <= r0[7];
cmp24_in1 <= r0[23];
r1[7] <= cmp24_out0;
r1[23] <= cmp24_out1;

cmp25_in0 <= r0[8];
cmp25_in1 <= r0[24];
r1[8] <= cmp25_out0;
r1[24] <= cmp25_out1;

cmp26_in0 <= r0[9];
cmp26_in1 <= r0[25];
r1[9] <= cmp26_out0;
r1[25] <= cmp26_out1;

cmp27_in0 <= r0[10];
cmp27_in1 <= r0[26];
r1[10] <= cmp27_out0;
r1[26] <= cmp27_out1;

cmp28_in0 <= r0[11];
cmp28_in1 <= r0[27];
r1[11] <= cmp28_out0;
r1[27] <= cmp28_out1;

cmp29_in0 <= r0[12];
cmp29_in1 <= r0[28];
r1[12] <= cmp29_out0;
r1[28] <= cmp29_out1;

cmp30_in0 <= r0[13];
cmp30_in1 <= r0[29];
r1[13] <= cmp30_out0;
r1[29] <= cmp30_out1;

cmp31_in0 <= r0[14];
cmp31_in1 <= r0[30];
r1[14] <= cmp31_out0;
r1[30] <= cmp31_out1;

cmp32_in0 <= r0[15];
cmp32_in1 <= r0[31];
r1[15] <= cmp32_out0;
r1[31] <= cmp32_out1;

cmp33_in0 <= r0[32];
cmp33_in1 <= r0[48];
r1[32] <= cmp33_out0;
r1[48] <= cmp33_out1;

r_1_33_tmp <= r0[33];
r1[33] <= r_1_33_tmp;

r_1_34_tmp <= r0[34];
r1[34] <= r_1_34_tmp;

r_1_35_tmp <= r0[35];
r1[35] <= r_1_35_tmp;

r_1_36_tmp <= r0[36];
r1[36] <= r_1_36_tmp;

r_1_37_tmp <= r0[37];
r1[37] <= r_1_37_tmp;

r_1_38_tmp <= r0[38];
r1[38] <= r_1_38_tmp;

r_1_39_tmp <= r0[39];
r1[39] <= r_1_39_tmp;

r_1_40_tmp <= r0[40];
r1[40] <= r_1_40_tmp;

r_1_41_tmp <= r0[41];
r1[41] <= r_1_41_tmp;

r_1_42_tmp <= r0[42];
r1[42] <= r_1_42_tmp;

r_1_43_tmp <= r0[43];
r1[43] <= r_1_43_tmp;

r_1_44_tmp <= r0[44];
r1[44] <= r_1_44_tmp;

r_1_45_tmp <= r0[45];
r1[45] <= r_1_45_tmp;

r_1_46_tmp <= r0[46];
r1[46] <= r_1_46_tmp;

r_1_47_tmp <= r0[47];
r1[47] <= r_1_47_tmp;

//--------------------------
//---------layer : 2------------
cmp34_in0 <= r1[16];
cmp34_in1 <= r1[32];
r2[16] <= cmp34_out0;
r2[32] <= cmp34_out1;

cmp35_in0 <= r1[17];
cmp35_in1 <= r1[33];
r2[17] <= cmp35_out0;
r2[33] <= cmp35_out1;

cmp36_in0 <= r1[18];
cmp36_in1 <= r1[34];
r2[18] <= cmp36_out0;
r2[34] <= cmp36_out1;

cmp37_in0 <= r1[19];
cmp37_in1 <= r1[35];
r2[19] <= cmp37_out0;
r2[35] <= cmp37_out1;

cmp38_in0 <= r1[20];
cmp38_in1 <= r1[36];
r2[20] <= cmp38_out0;
r2[36] <= cmp38_out1;

cmp39_in0 <= r1[21];
cmp39_in1 <= r1[37];
r2[21] <= cmp39_out0;
r2[37] <= cmp39_out1;

cmp40_in0 <= r1[22];
cmp40_in1 <= r1[38];
r2[22] <= cmp40_out0;
r2[38] <= cmp40_out1;

cmp41_in0 <= r1[23];
cmp41_in1 <= r1[39];
r2[23] <= cmp41_out0;
r2[39] <= cmp41_out1;

cmp42_in0 <= r1[24];
cmp42_in1 <= r1[40];
r2[24] <= cmp42_out0;
r2[40] <= cmp42_out1;

cmp43_in0 <= r1[25];
cmp43_in1 <= r1[41];
r2[25] <= cmp43_out0;
r2[41] <= cmp43_out1;

cmp44_in0 <= r1[26];
cmp44_in1 <= r1[42];
r2[26] <= cmp44_out0;
r2[42] <= cmp44_out1;

cmp45_in0 <= r1[27];
cmp45_in1 <= r1[43];
r2[27] <= cmp45_out0;
r2[43] <= cmp45_out1;

cmp46_in0 <= r1[28];
cmp46_in1 <= r1[44];
r2[28] <= cmp46_out0;
r2[44] <= cmp46_out1;

cmp47_in0 <= r1[29];
cmp47_in1 <= r1[45];
r2[29] <= cmp47_out0;
r2[45] <= cmp47_out1;

cmp48_in0 <= r1[30];
cmp48_in1 <= r1[46];
r2[30] <= cmp48_out0;
r2[46] <= cmp48_out1;

cmp49_in0 <= r1[31];
cmp49_in1 <= r1[47];
r2[31] <= cmp49_out0;
r2[47] <= cmp49_out1;

cmp50_in0 <= r1[0];
cmp50_in1 <= r1[8];
r2[0] <= cmp50_out0;
r2[8] <= cmp50_out1;

cmp51_in0 <= r1[1];
cmp51_in1 <= r1[9];
r2[1] <= cmp51_out0;
r2[9] <= cmp51_out1;

cmp52_in0 <= r1[2];
cmp52_in1 <= r1[10];
r2[2] <= cmp52_out0;
r2[10] <= cmp52_out1;

cmp53_in0 <= r1[3];
cmp53_in1 <= r1[11];
r2[3] <= cmp53_out0;
r2[11] <= cmp53_out1;

cmp54_in0 <= r1[4];
cmp54_in1 <= r1[12];
r2[4] <= cmp54_out0;
r2[12] <= cmp54_out1;

cmp55_in0 <= r1[5];
cmp55_in1 <= r1[13];
r2[5] <= cmp55_out0;
r2[13] <= cmp55_out1;

cmp56_in0 <= r1[6];
cmp56_in1 <= r1[14];
r2[6] <= cmp56_out0;
r2[14] <= cmp56_out1;

cmp57_in0 <= r1[7];
cmp57_in1 <= r1[15];
r2[7] <= cmp57_out0;
r2[15] <= cmp57_out1;

r_2_48_tmp <= r1[48];
r2[48] <= r_2_48_tmp;

//--------------------------
//---------layer : 3------------
cmp58_in0 <= r2[16];
cmp58_in1 <= r2[24];
r3[16] <= cmp58_out0;
r3[24] <= cmp58_out1;

cmp59_in0 <= r2[17];
cmp59_in1 <= r2[25];
r3[17] <= cmp59_out0;
r3[25] <= cmp59_out1;

cmp60_in0 <= r2[18];
cmp60_in1 <= r2[26];
r3[18] <= cmp60_out0;
r3[26] <= cmp60_out1;

cmp61_in0 <= r2[19];
cmp61_in1 <= r2[27];
r3[19] <= cmp61_out0;
r3[27] <= cmp61_out1;

cmp62_in0 <= r2[20];
cmp62_in1 <= r2[28];
r3[20] <= cmp62_out0;
r3[28] <= cmp62_out1;

cmp63_in0 <= r2[21];
cmp63_in1 <= r2[29];
r3[21] <= cmp63_out0;
r3[29] <= cmp63_out1;

cmp64_in0 <= r2[22];
cmp64_in1 <= r2[30];
r3[22] <= cmp64_out0;
r3[30] <= cmp64_out1;

cmp65_in0 <= r2[23];
cmp65_in1 <= r2[31];
r3[23] <= cmp65_out0;
r3[31] <= cmp65_out1;

cmp66_in0 <= r2[32];
cmp66_in1 <= r2[40];
r3[32] <= cmp66_out0;
r3[40] <= cmp66_out1;

cmp67_in0 <= r2[33];
cmp67_in1 <= r2[41];
r3[33] <= cmp67_out0;
r3[41] <= cmp67_out1;

cmp68_in0 <= r2[34];
cmp68_in1 <= r2[42];
r3[34] <= cmp68_out0;
r3[42] <= cmp68_out1;

cmp69_in0 <= r2[35];
cmp69_in1 <= r2[43];
r3[35] <= cmp69_out0;
r3[43] <= cmp69_out1;

cmp70_in0 <= r2[36];
cmp70_in1 <= r2[44];
r3[36] <= cmp70_out0;
r3[44] <= cmp70_out1;

cmp71_in0 <= r2[37];
cmp71_in1 <= r2[45];
r3[37] <= cmp71_out0;
r3[45] <= cmp71_out1;

cmp72_in0 <= r2[38];
cmp72_in1 <= r2[46];
r3[38] <= cmp72_out0;
r3[46] <= cmp72_out1;

cmp73_in0 <= r2[39];
cmp73_in1 <= r2[47];
r3[39] <= cmp73_out0;
r3[47] <= cmp73_out1;

r_3_0_tmp <= r2[0];
r3[0] <= r_3_0_tmp;

r_3_1_tmp <= r2[1];
r3[1] <= r_3_1_tmp;

r_3_2_tmp <= r2[2];
r3[2] <= r_3_2_tmp;

r_3_3_tmp <= r2[3];
r3[3] <= r_3_3_tmp;

r_3_4_tmp <= r2[4];
r3[4] <= r_3_4_tmp;

r_3_5_tmp <= r2[5];
r3[5] <= r_3_5_tmp;

r_3_6_tmp <= r2[6];
r3[6] <= r_3_6_tmp;

r_3_7_tmp <= r2[7];
r3[7] <= r_3_7_tmp;

r_3_8_tmp <= r2[8];
r3[8] <= r_3_8_tmp;

r_3_9_tmp <= r2[9];
r3[9] <= r_3_9_tmp;

r_3_10_tmp <= r2[10];
r3[10] <= r_3_10_tmp;

r_3_11_tmp <= r2[11];
r3[11] <= r_3_11_tmp;

r_3_12_tmp <= r2[12];
r3[12] <= r_3_12_tmp;

r_3_13_tmp <= r2[13];
r3[13] <= r_3_13_tmp;

r_3_14_tmp <= r2[14];
r3[14] <= r_3_14_tmp;

r_3_15_tmp <= r2[15];
r3[15] <= r_3_15_tmp;

r_3_48_tmp <= r2[48];
r3[48] <= r_3_48_tmp;

//--------------------------
//---------layer : 4------------
cmp74_in0 <= r3[8];
cmp74_in1 <= r3[32];
r4[8] <= cmp74_out0;
r4[32] <= cmp74_out1;

cmp75_in0 <= r3[9];
cmp75_in1 <= r3[33];
r4[9] <= cmp75_out0;
r4[33] <= cmp75_out1;

cmp76_in0 <= r3[10];
cmp76_in1 <= r3[34];
r4[10] <= cmp76_out0;
r4[34] <= cmp76_out1;

cmp77_in0 <= r3[11];
cmp77_in1 <= r3[35];
r4[11] <= cmp77_out0;
r4[35] <= cmp77_out1;

cmp78_in0 <= r3[12];
cmp78_in1 <= r3[36];
r4[12] <= cmp78_out0;
r4[36] <= cmp78_out1;

cmp79_in0 <= r3[13];
cmp79_in1 <= r3[37];
r4[13] <= cmp79_out0;
r4[37] <= cmp79_out1;

cmp80_in0 <= r3[14];
cmp80_in1 <= r3[38];
r4[14] <= cmp80_out0;
r4[38] <= cmp80_out1;

cmp81_in0 <= r3[15];
cmp81_in1 <= r3[39];
r4[15] <= cmp81_out0;
r4[39] <= cmp81_out1;

cmp82_in0 <= r3[24];
cmp82_in1 <= r3[48];
r4[24] <= cmp82_out0;
r4[48] <= cmp82_out1;

r_4_0_tmp <= r3[0];
r4[0] <= r_4_0_tmp;

r_4_1_tmp <= r3[1];
r4[1] <= r_4_1_tmp;

r_4_2_tmp <= r3[2];
r4[2] <= r_4_2_tmp;

r_4_3_tmp <= r3[3];
r4[3] <= r_4_3_tmp;

r_4_4_tmp <= r3[4];
r4[4] <= r_4_4_tmp;

r_4_5_tmp <= r3[5];
r4[5] <= r_4_5_tmp;

r_4_6_tmp <= r3[6];
r4[6] <= r_4_6_tmp;

r_4_7_tmp <= r3[7];
r4[7] <= r_4_7_tmp;

r_4_16_tmp <= r3[16];
r4[16] <= r_4_16_tmp;

r_4_17_tmp <= r3[17];
r4[17] <= r_4_17_tmp;

r_4_18_tmp <= r3[18];
r4[18] <= r_4_18_tmp;

r_4_19_tmp <= r3[19];
r4[19] <= r_4_19_tmp;

r_4_20_tmp <= r3[20];
r4[20] <= r_4_20_tmp;

r_4_21_tmp <= r3[21];
r4[21] <= r_4_21_tmp;

r_4_22_tmp <= r3[22];
r4[22] <= r_4_22_tmp;

r_4_23_tmp <= r3[23];
r4[23] <= r_4_23_tmp;

r_4_25_tmp <= r3[25];
r4[25] <= r_4_25_tmp;

r_4_26_tmp <= r3[26];
r4[26] <= r_4_26_tmp;

r_4_27_tmp <= r3[27];
r4[27] <= r_4_27_tmp;

r_4_28_tmp <= r3[28];
r4[28] <= r_4_28_tmp;

r_4_29_tmp <= r3[29];
r4[29] <= r_4_29_tmp;

r_4_30_tmp <= r3[30];
r4[30] <= r_4_30_tmp;

r_4_31_tmp <= r3[31];
r4[31] <= r_4_31_tmp;

r_4_40_tmp <= r3[40];
r4[40] <= r_4_40_tmp;

r_4_41_tmp <= r3[41];
r4[41] <= r_4_41_tmp;

r_4_42_tmp <= r3[42];
r4[42] <= r_4_42_tmp;

r_4_43_tmp <= r3[43];
r4[43] <= r_4_43_tmp;

r_4_44_tmp <= r3[44];
r4[44] <= r_4_44_tmp;

r_4_45_tmp <= r3[45];
r4[45] <= r_4_45_tmp;

r_4_46_tmp <= r3[46];
r4[46] <= r_4_46_tmp;

r_4_47_tmp <= r3[47];
r4[47] <= r_4_47_tmp;

//--------------------------
//---------layer : 5------------
cmp83_in0 <= r4[8];
cmp83_in1 <= r4[16];
r5[8] <= cmp83_out0;
r5[16] <= cmp83_out1;

cmp84_in0 <= r4[9];
cmp84_in1 <= r4[17];
r5[9] <= cmp84_out0;
r5[17] <= cmp84_out1;

cmp85_in0 <= r4[10];
cmp85_in1 <= r4[18];
r5[10] <= cmp85_out0;
r5[18] <= cmp85_out1;

cmp86_in0 <= r4[11];
cmp86_in1 <= r4[19];
r5[11] <= cmp86_out0;
r5[19] <= cmp86_out1;

cmp87_in0 <= r4[12];
cmp87_in1 <= r4[20];
r5[12] <= cmp87_out0;
r5[20] <= cmp87_out1;

cmp88_in0 <= r4[13];
cmp88_in1 <= r4[21];
r5[13] <= cmp88_out0;
r5[21] <= cmp88_out1;

cmp89_in0 <= r4[14];
cmp89_in1 <= r4[22];
r5[14] <= cmp89_out0;
r5[22] <= cmp89_out1;

cmp90_in0 <= r4[15];
cmp90_in1 <= r4[23];
r5[15] <= cmp90_out0;
r5[23] <= cmp90_out1;

cmp91_in0 <= r4[24];
cmp91_in1 <= r4[32];
r5[24] <= cmp91_out0;
r5[32] <= cmp91_out1;

cmp92_in0 <= r4[25];
cmp92_in1 <= r4[33];
r5[25] <= cmp92_out0;
r5[33] <= cmp92_out1;

cmp93_in0 <= r4[26];
cmp93_in1 <= r4[34];
r5[26] <= cmp93_out0;
r5[34] <= cmp93_out1;

cmp94_in0 <= r4[27];
cmp94_in1 <= r4[35];
r5[27] <= cmp94_out0;
r5[35] <= cmp94_out1;

cmp95_in0 <= r4[28];
cmp95_in1 <= r4[36];
r5[28] <= cmp95_out0;
r5[36] <= cmp95_out1;

cmp96_in0 <= r4[29];
cmp96_in1 <= r4[37];
r5[29] <= cmp96_out0;
r5[37] <= cmp96_out1;

cmp97_in0 <= r4[30];
cmp97_in1 <= r4[38];
r5[30] <= cmp97_out0;
r5[38] <= cmp97_out1;

cmp98_in0 <= r4[31];
cmp98_in1 <= r4[39];
r5[31] <= cmp98_out0;
r5[39] <= cmp98_out1;

cmp99_in0 <= r4[40];
cmp99_in1 <= r4[48];
r5[40] <= cmp99_out0;
r5[48] <= cmp99_out1;

cmp100_in0 <= r4[0];
cmp100_in1 <= r4[4];
r5[0] <= cmp100_out0;
r5[4] <= cmp100_out1;

cmp101_in0 <= r4[1];
cmp101_in1 <= r4[5];
r5[1] <= cmp101_out0;
r5[5] <= cmp101_out1;

cmp102_in0 <= r4[2];
cmp102_in1 <= r4[6];
r5[2] <= cmp102_out0;
r5[6] <= cmp102_out1;

cmp103_in0 <= r4[3];
cmp103_in1 <= r4[7];
r5[3] <= cmp103_out0;
r5[7] <= cmp103_out1;

r_5_41_tmp <= r4[41];
r5[41] <= r_5_41_tmp;

r_5_42_tmp <= r4[42];
r5[42] <= r_5_42_tmp;

r_5_43_tmp <= r4[43];
r5[43] <= r_5_43_tmp;

r_5_44_tmp <= r4[44];
r5[44] <= r_5_44_tmp;

r_5_45_tmp <= r4[45];
r5[45] <= r_5_45_tmp;

r_5_46_tmp <= r4[46];
r5[46] <= r_5_46_tmp;

r_5_47_tmp <= r4[47];
r5[47] <= r_5_47_tmp;

//--------------------------
//---------layer : 6------------
cmp104_in0 <= r5[8];
cmp104_in1 <= r5[12];
r6[8] <= cmp104_out0;
r6[12] <= cmp104_out1;

cmp105_in0 <= r5[9];
cmp105_in1 <= r5[13];
r6[9] <= cmp105_out0;
r6[13] <= cmp105_out1;

cmp106_in0 <= r5[10];
cmp106_in1 <= r5[14];
r6[10] <= cmp106_out0;
r6[14] <= cmp106_out1;

cmp107_in0 <= r5[11];
cmp107_in1 <= r5[15];
r6[11] <= cmp107_out0;
r6[15] <= cmp107_out1;

cmp108_in0 <= r5[16];
cmp108_in1 <= r5[20];
r6[16] <= cmp108_out0;
r6[20] <= cmp108_out1;

cmp109_in0 <= r5[17];
cmp109_in1 <= r5[21];
r6[17] <= cmp109_out0;
r6[21] <= cmp109_out1;

cmp110_in0 <= r5[18];
cmp110_in1 <= r5[22];
r6[18] <= cmp110_out0;
r6[22] <= cmp110_out1;

cmp111_in0 <= r5[19];
cmp111_in1 <= r5[23];
r6[19] <= cmp111_out0;
r6[23] <= cmp111_out1;

cmp112_in0 <= r5[24];
cmp112_in1 <= r5[28];
r6[24] <= cmp112_out0;
r6[28] <= cmp112_out1;

cmp113_in0 <= r5[25];
cmp113_in1 <= r5[29];
r6[25] <= cmp113_out0;
r6[29] <= cmp113_out1;

cmp114_in0 <= r5[26];
cmp114_in1 <= r5[30];
r6[26] <= cmp114_out0;
r6[30] <= cmp114_out1;

cmp115_in0 <= r5[27];
cmp115_in1 <= r5[31];
r6[27] <= cmp115_out0;
r6[31] <= cmp115_out1;

cmp116_in0 <= r5[32];
cmp116_in1 <= r5[36];
r6[32] <= cmp116_out0;
r6[36] <= cmp116_out1;

cmp117_in0 <= r5[33];
cmp117_in1 <= r5[37];
r6[33] <= cmp117_out0;
r6[37] <= cmp117_out1;

cmp118_in0 <= r5[34];
cmp118_in1 <= r5[38];
r6[34] <= cmp118_out0;
r6[38] <= cmp118_out1;

cmp119_in0 <= r5[35];
cmp119_in1 <= r5[39];
r6[35] <= cmp119_out0;
r6[39] <= cmp119_out1;

cmp120_in0 <= r5[40];
cmp120_in1 <= r5[44];
r6[40] <= cmp120_out0;
r6[44] <= cmp120_out1;

cmp121_in0 <= r5[41];
cmp121_in1 <= r5[45];
r6[41] <= cmp121_out0;
r6[45] <= cmp121_out1;

cmp122_in0 <= r5[42];
cmp122_in1 <= r5[46];
r6[42] <= cmp122_out0;
r6[46] <= cmp122_out1;

cmp123_in0 <= r5[43];
cmp123_in1 <= r5[47];
r6[43] <= cmp123_out0;
r6[47] <= cmp123_out1;

r_6_0_tmp <= r5[0];
r6[0] <= r_6_0_tmp;

r_6_1_tmp <= r5[1];
r6[1] <= r_6_1_tmp;

r_6_2_tmp <= r5[2];
r6[2] <= r_6_2_tmp;

r_6_3_tmp <= r5[3];
r6[3] <= r_6_3_tmp;

r_6_4_tmp <= r5[4];
r6[4] <= r_6_4_tmp;

r_6_5_tmp <= r5[5];
r6[5] <= r_6_5_tmp;

r_6_6_tmp <= r5[6];
r6[6] <= r_6_6_tmp;

r_6_7_tmp <= r5[7];
r6[7] <= r_6_7_tmp;

r_6_48_tmp <= r5[48];
r6[48] <= r_6_48_tmp;

//--------------------------
//---------layer : 7------------
cmp124_in0 <= r6[4];
cmp124_in1 <= r6[32];
r7[4] <= cmp124_out0;
r7[32] <= cmp124_out1;

cmp125_in0 <= r6[5];
cmp125_in1 <= r6[33];
r7[5] <= cmp125_out0;
r7[33] <= cmp125_out1;

cmp126_in0 <= r6[6];
cmp126_in1 <= r6[34];
r7[6] <= cmp126_out0;
r7[34] <= cmp126_out1;

cmp127_in0 <= r6[7];
cmp127_in1 <= r6[35];
r7[7] <= cmp127_out0;
r7[35] <= cmp127_out1;

cmp128_in0 <= r6[12];
cmp128_in1 <= r6[40];
r7[12] <= cmp128_out0;
r7[40] <= cmp128_out1;

cmp129_in0 <= r6[13];
cmp129_in1 <= r6[41];
r7[13] <= cmp129_out0;
r7[41] <= cmp129_out1;

cmp130_in0 <= r6[14];
cmp130_in1 <= r6[42];
r7[14] <= cmp130_out0;
r7[42] <= cmp130_out1;

cmp131_in0 <= r6[15];
cmp131_in1 <= r6[43];
r7[15] <= cmp131_out0;
r7[43] <= cmp131_out1;

cmp132_in0 <= r6[20];
cmp132_in1 <= r6[48];
r7[20] <= cmp132_out0;
r7[48] <= cmp132_out1;

r_7_0_tmp <= r6[0];
r7[0] <= r_7_0_tmp;

r_7_1_tmp <= r6[1];
r7[1] <= r_7_1_tmp;

r_7_2_tmp <= r6[2];
r7[2] <= r_7_2_tmp;

r_7_3_tmp <= r6[3];
r7[3] <= r_7_3_tmp;

r_7_8_tmp <= r6[8];
r7[8] <= r_7_8_tmp;

r_7_9_tmp <= r6[9];
r7[9] <= r_7_9_tmp;

r_7_10_tmp <= r6[10];
r7[10] <= r_7_10_tmp;

r_7_11_tmp <= r6[11];
r7[11] <= r_7_11_tmp;

r_7_16_tmp <= r6[16];
r7[16] <= r_7_16_tmp;

r_7_17_tmp <= r6[17];
r7[17] <= r_7_17_tmp;

r_7_18_tmp <= r6[18];
r7[18] <= r_7_18_tmp;

r_7_19_tmp <= r6[19];
r7[19] <= r_7_19_tmp;

r_7_21_tmp <= r6[21];
r7[21] <= r_7_21_tmp;

r_7_22_tmp <= r6[22];
r7[22] <= r_7_22_tmp;

r_7_23_tmp <= r6[23];
r7[23] <= r_7_23_tmp;

r_7_24_tmp <= r6[24];
r7[24] <= r_7_24_tmp;

r_7_25_tmp <= r6[25];
r7[25] <= r_7_25_tmp;

r_7_26_tmp <= r6[26];
r7[26] <= r_7_26_tmp;

r_7_27_tmp <= r6[27];
r7[27] <= r_7_27_tmp;

r_7_28_tmp <= r6[28];
r7[28] <= r_7_28_tmp;

r_7_29_tmp <= r6[29];
r7[29] <= r_7_29_tmp;

r_7_30_tmp <= r6[30];
r7[30] <= r_7_30_tmp;

r_7_31_tmp <= r6[31];
r7[31] <= r_7_31_tmp;

r_7_36_tmp <= r6[36];
r7[36] <= r_7_36_tmp;

r_7_37_tmp <= r6[37];
r7[37] <= r_7_37_tmp;

r_7_38_tmp <= r6[38];
r7[38] <= r_7_38_tmp;

r_7_39_tmp <= r6[39];
r7[39] <= r_7_39_tmp;

r_7_44_tmp <= r6[44];
r7[44] <= r_7_44_tmp;

r_7_45_tmp <= r6[45];
r7[45] <= r_7_45_tmp;

r_7_46_tmp <= r6[46];
r7[46] <= r_7_46_tmp;

r_7_47_tmp <= r6[47];
r7[47] <= r_7_47_tmp;

//--------------------------
//---------layer : 8------------
cmp133_in0 <= r7[4];
cmp133_in1 <= r7[16];
r8[4] <= cmp133_out0;
r8[16] <= cmp133_out1;

cmp134_in0 <= r7[5];
cmp134_in1 <= r7[17];
r8[5] <= cmp134_out0;
r8[17] <= cmp134_out1;

cmp135_in0 <= r7[6];
cmp135_in1 <= r7[18];
r8[6] <= cmp135_out0;
r8[18] <= cmp135_out1;

cmp136_in0 <= r7[7];
cmp136_in1 <= r7[19];
r8[7] <= cmp136_out0;
r8[19] <= cmp136_out1;

cmp137_in0 <= r7[12];
cmp137_in1 <= r7[24];
r8[12] <= cmp137_out0;
r8[24] <= cmp137_out1;

cmp138_in0 <= r7[13];
cmp138_in1 <= r7[25];
r8[13] <= cmp138_out0;
r8[25] <= cmp138_out1;

cmp139_in0 <= r7[14];
cmp139_in1 <= r7[26];
r8[14] <= cmp139_out0;
r8[26] <= cmp139_out1;

cmp140_in0 <= r7[15];
cmp140_in1 <= r7[27];
r8[15] <= cmp140_out0;
r8[27] <= cmp140_out1;

cmp141_in0 <= r7[20];
cmp141_in1 <= r7[32];
r8[20] <= cmp141_out0;
r8[32] <= cmp141_out1;

cmp142_in0 <= r7[21];
cmp142_in1 <= r7[33];
r8[21] <= cmp142_out0;
r8[33] <= cmp142_out1;

cmp143_in0 <= r7[22];
cmp143_in1 <= r7[34];
r8[22] <= cmp143_out0;
r8[34] <= cmp143_out1;

cmp144_in0 <= r7[23];
cmp144_in1 <= r7[35];
r8[23] <= cmp144_out0;
r8[35] <= cmp144_out1;

cmp145_in0 <= r7[28];
cmp145_in1 <= r7[40];
r8[28] <= cmp145_out0;
r8[40] <= cmp145_out1;

cmp146_in0 <= r7[29];
cmp146_in1 <= r7[41];
r8[29] <= cmp146_out0;
r8[41] <= cmp146_out1;

cmp147_in0 <= r7[30];
cmp147_in1 <= r7[42];
r8[30] <= cmp147_out0;
r8[42] <= cmp147_out1;

cmp148_in0 <= r7[31];
cmp148_in1 <= r7[43];
r8[31] <= cmp148_out0;
r8[43] <= cmp148_out1;

cmp149_in0 <= r7[36];
cmp149_in1 <= r7[48];
r8[36] <= cmp149_out0;
r8[48] <= cmp149_out1;

r_8_0_tmp <= r7[0];
r8[0] <= r_8_0_tmp;

r_8_1_tmp <= r7[1];
r8[1] <= r_8_1_tmp;

r_8_2_tmp <= r7[2];
r8[2] <= r_8_2_tmp;

r_8_3_tmp <= r7[3];
r8[3] <= r_8_3_tmp;

r_8_8_tmp <= r7[8];
r8[8] <= r_8_8_tmp;

r_8_9_tmp <= r7[9];
r8[9] <= r_8_9_tmp;

r_8_10_tmp <= r7[10];
r8[10] <= r_8_10_tmp;

r_8_11_tmp <= r7[11];
r8[11] <= r_8_11_tmp;

r_8_37_tmp <= r7[37];
r8[37] <= r_8_37_tmp;

r_8_38_tmp <= r7[38];
r8[38] <= r_8_38_tmp;

r_8_39_tmp <= r7[39];
r8[39] <= r_8_39_tmp;

r_8_44_tmp <= r7[44];
r8[44] <= r_8_44_tmp;

r_8_45_tmp <= r7[45];
r8[45] <= r_8_45_tmp;

r_8_46_tmp <= r7[46];
r8[46] <= r_8_46_tmp;

r_8_47_tmp <= r7[47];
r8[47] <= r_8_47_tmp;

//--------------------------
//---------layer : 9------------
cmp150_in0 <= r8[4];
cmp150_in1 <= r8[8];
r9[4] <= cmp150_out0;
r9[8] <= cmp150_out1;

cmp151_in0 <= r8[5];
cmp151_in1 <= r8[9];
r9[5] <= cmp151_out0;
r9[9] <= cmp151_out1;

cmp152_in0 <= r8[6];
cmp152_in1 <= r8[10];
r9[6] <= cmp152_out0;
r9[10] <= cmp152_out1;

cmp153_in0 <= r8[7];
cmp153_in1 <= r8[11];
r9[7] <= cmp153_out0;
r9[11] <= cmp153_out1;

cmp154_in0 <= r8[12];
cmp154_in1 <= r8[16];
r9[12] <= cmp154_out0;
r9[16] <= cmp154_out1;

cmp155_in0 <= r8[13];
cmp155_in1 <= r8[17];
r9[13] <= cmp155_out0;
r9[17] <= cmp155_out1;

cmp156_in0 <= r8[14];
cmp156_in1 <= r8[18];
r9[14] <= cmp156_out0;
r9[18] <= cmp156_out1;

cmp157_in0 <= r8[15];
cmp157_in1 <= r8[19];
r9[15] <= cmp157_out0;
r9[19] <= cmp157_out1;

cmp158_in0 <= r8[20];
cmp158_in1 <= r8[24];
r9[20] <= cmp158_out0;
r9[24] <= cmp158_out1;

cmp159_in0 <= r8[21];
cmp159_in1 <= r8[25];
r9[21] <= cmp159_out0;
r9[25] <= cmp159_out1;

cmp160_in0 <= r8[22];
cmp160_in1 <= r8[26];
r9[22] <= cmp160_out0;
r9[26] <= cmp160_out1;

cmp161_in0 <= r8[23];
cmp161_in1 <= r8[27];
r9[23] <= cmp161_out0;
r9[27] <= cmp161_out1;

cmp162_in0 <= r8[28];
cmp162_in1 <= r8[32];
r9[28] <= cmp162_out0;
r9[32] <= cmp162_out1;

cmp163_in0 <= r8[29];
cmp163_in1 <= r8[33];
r9[29] <= cmp163_out0;
r9[33] <= cmp163_out1;

cmp164_in0 <= r8[30];
cmp164_in1 <= r8[34];
r9[30] <= cmp164_out0;
r9[34] <= cmp164_out1;

cmp165_in0 <= r8[31];
cmp165_in1 <= r8[35];
r9[31] <= cmp165_out0;
r9[35] <= cmp165_out1;

cmp166_in0 <= r8[36];
cmp166_in1 <= r8[40];
r9[36] <= cmp166_out0;
r9[40] <= cmp166_out1;

cmp167_in0 <= r8[37];
cmp167_in1 <= r8[41];
r9[37] <= cmp167_out0;
r9[41] <= cmp167_out1;

cmp168_in0 <= r8[38];
cmp168_in1 <= r8[42];
r9[38] <= cmp168_out0;
r9[42] <= cmp168_out1;

cmp169_in0 <= r8[39];
cmp169_in1 <= r8[43];
r9[39] <= cmp169_out0;
r9[43] <= cmp169_out1;

cmp170_in0 <= r8[44];
cmp170_in1 <= r8[48];
r9[44] <= cmp170_out0;
r9[48] <= cmp170_out1;

cmp171_in0 <= r8[0];
cmp171_in1 <= r8[2];
r9[0] <= cmp171_out0;
r9[2] <= cmp171_out1;

cmp172_in0 <= r8[1];
cmp172_in1 <= r8[3];
r9[1] <= cmp172_out0;
r9[3] <= cmp172_out1;

r_9_45_tmp <= r8[45];
r9[45] <= r_9_45_tmp;

r_9_46_tmp <= r8[46];
r9[46] <= r_9_46_tmp;

r_9_47_tmp <= r8[47];
r9[47] <= r_9_47_tmp;

//--------------------------
//---------layer : 10------------
cmp173_in0 <= r9[4];
cmp173_in1 <= r9[6];
r10[4] <= cmp173_out0;
r10[6] <= cmp173_out1;

cmp174_in0 <= r9[5];
cmp174_in1 <= r9[7];
r10[5] <= cmp174_out0;
r10[7] <= cmp174_out1;

cmp175_in0 <= r9[8];
cmp175_in1 <= r9[10];
r10[8] <= cmp175_out0;
r10[10] <= cmp175_out1;

cmp176_in0 <= r9[9];
cmp176_in1 <= r9[11];
r10[9] <= cmp176_out0;
r10[11] <= cmp176_out1;

cmp177_in0 <= r9[12];
cmp177_in1 <= r9[14];
r10[12] <= cmp177_out0;
r10[14] <= cmp177_out1;

cmp178_in0 <= r9[13];
cmp178_in1 <= r9[15];
r10[13] <= cmp178_out0;
r10[15] <= cmp178_out1;

cmp179_in0 <= r9[16];
cmp179_in1 <= r9[18];
r10[16] <= cmp179_out0;
r10[18] <= cmp179_out1;

cmp180_in0 <= r9[17];
cmp180_in1 <= r9[19];
r10[17] <= cmp180_out0;
r10[19] <= cmp180_out1;

cmp181_in0 <= r9[20];
cmp181_in1 <= r9[22];
r10[20] <= cmp181_out0;
r10[22] <= cmp181_out1;

cmp182_in0 <= r9[21];
cmp182_in1 <= r9[23];
r10[21] <= cmp182_out0;
r10[23] <= cmp182_out1;

cmp183_in0 <= r9[24];
cmp183_in1 <= r9[26];
r10[24] <= cmp183_out0;
r10[26] <= cmp183_out1;

cmp184_in0 <= r9[25];
cmp184_in1 <= r9[27];
r10[25] <= cmp184_out0;
r10[27] <= cmp184_out1;

cmp185_in0 <= r9[28];
cmp185_in1 <= r9[30];
r10[28] <= cmp185_out0;
r10[30] <= cmp185_out1;

cmp186_in0 <= r9[29];
cmp186_in1 <= r9[31];
r10[29] <= cmp186_out0;
r10[31] <= cmp186_out1;

cmp187_in0 <= r9[32];
cmp187_in1 <= r9[34];
r10[32] <= cmp187_out0;
r10[34] <= cmp187_out1;

cmp188_in0 <= r9[33];
cmp188_in1 <= r9[35];
r10[33] <= cmp188_out0;
r10[35] <= cmp188_out1;

cmp189_in0 <= r9[36];
cmp189_in1 <= r9[38];
r10[36] <= cmp189_out0;
r10[38] <= cmp189_out1;

cmp190_in0 <= r9[37];
cmp190_in1 <= r9[39];
r10[37] <= cmp190_out0;
r10[39] <= cmp190_out1;

cmp191_in0 <= r9[40];
cmp191_in1 <= r9[42];
r10[40] <= cmp191_out0;
r10[42] <= cmp191_out1;

cmp192_in0 <= r9[41];
cmp192_in1 <= r9[43];
r10[41] <= cmp192_out0;
r10[43] <= cmp192_out1;

cmp193_in0 <= r9[44];
cmp193_in1 <= r9[46];
r10[44] <= cmp193_out0;
r10[46] <= cmp193_out1;

cmp194_in0 <= r9[45];
cmp194_in1 <= r9[47];
r10[45] <= cmp194_out0;
r10[47] <= cmp194_out1;

r_10_0_tmp <= r9[0];
r10[0] <= r_10_0_tmp;

r_10_1_tmp <= r9[1];
r10[1] <= r_10_1_tmp;

r_10_2_tmp <= r9[2];
r10[2] <= r_10_2_tmp;

r_10_3_tmp <= r9[3];
r10[3] <= r_10_3_tmp;

r_10_48_tmp <= r9[48];
r10[48] <= r_10_48_tmp;

//--------------------------
//---------layer : 11------------
cmp195_in0 <= r10[2];
cmp195_in1 <= r10[32];
r11[2] <= cmp195_out0;
r11[32] <= cmp195_out1;

cmp196_in0 <= r10[3];
cmp196_in1 <= r10[33];
r11[3] <= cmp196_out0;
r11[33] <= cmp196_out1;

cmp197_in0 <= r10[6];
cmp197_in1 <= r10[36];
r11[6] <= cmp197_out0;
r11[36] <= cmp197_out1;

cmp198_in0 <= r10[7];
cmp198_in1 <= r10[37];
r11[7] <= cmp198_out0;
r11[37] <= cmp198_out1;

cmp199_in0 <= r10[10];
cmp199_in1 <= r10[40];
r11[10] <= cmp199_out0;
r11[40] <= cmp199_out1;

cmp200_in0 <= r10[11];
cmp200_in1 <= r10[41];
r11[11] <= cmp200_out0;
r11[41] <= cmp200_out1;

cmp201_in0 <= r10[14];
cmp201_in1 <= r10[44];
r11[14] <= cmp201_out0;
r11[44] <= cmp201_out1;

cmp202_in0 <= r10[15];
cmp202_in1 <= r10[45];
r11[15] <= cmp202_out0;
r11[45] <= cmp202_out1;

cmp203_in0 <= r10[18];
cmp203_in1 <= r10[48];
r11[18] <= cmp203_out0;
r11[48] <= cmp203_out1;

r_11_0_tmp <= r10[0];
r11[0] <= r_11_0_tmp;

r_11_1_tmp <= r10[1];
r11[1] <= r_11_1_tmp;

r_11_4_tmp <= r10[4];
r11[4] <= r_11_4_tmp;

r_11_5_tmp <= r10[5];
r11[5] <= r_11_5_tmp;

r_11_8_tmp <= r10[8];
r11[8] <= r_11_8_tmp;

r_11_9_tmp <= r10[9];
r11[9] <= r_11_9_tmp;

r_11_12_tmp <= r10[12];
r11[12] <= r_11_12_tmp;

r_11_13_tmp <= r10[13];
r11[13] <= r_11_13_tmp;

r_11_16_tmp <= r10[16];
r11[16] <= r_11_16_tmp;

r_11_17_tmp <= r10[17];
r11[17] <= r_11_17_tmp;

r_11_19_tmp <= r10[19];
r11[19] <= r_11_19_tmp;

r_11_20_tmp <= r10[20];
r11[20] <= r_11_20_tmp;

r_11_21_tmp <= r10[21];
r11[21] <= r_11_21_tmp;

r_11_22_tmp <= r10[22];
r11[22] <= r_11_22_tmp;

r_11_23_tmp <= r10[23];
r11[23] <= r_11_23_tmp;

r_11_24_tmp <= r10[24];
r11[24] <= r_11_24_tmp;

r_11_25_tmp <= r10[25];
r11[25] <= r_11_25_tmp;

r_11_26_tmp <= r10[26];
r11[26] <= r_11_26_tmp;

r_11_27_tmp <= r10[27];
r11[27] <= r_11_27_tmp;

r_11_28_tmp <= r10[28];
r11[28] <= r_11_28_tmp;

r_11_29_tmp <= r10[29];
r11[29] <= r_11_29_tmp;

r_11_30_tmp <= r10[30];
r11[30] <= r_11_30_tmp;

r_11_31_tmp <= r10[31];
r11[31] <= r_11_31_tmp;

r_11_34_tmp <= r10[34];
r11[34] <= r_11_34_tmp;

r_11_35_tmp <= r10[35];
r11[35] <= r_11_35_tmp;

r_11_38_tmp <= r10[38];
r11[38] <= r_11_38_tmp;

r_11_39_tmp <= r10[39];
r11[39] <= r_11_39_tmp;

r_11_42_tmp <= r10[42];
r11[42] <= r_11_42_tmp;

r_11_43_tmp <= r10[43];
r11[43] <= r_11_43_tmp;

r_11_46_tmp <= r10[46];
r11[46] <= r_11_46_tmp;

r_11_47_tmp <= r10[47];
r11[47] <= r_11_47_tmp;

//--------------------------
//---------layer : 12------------
cmp204_in0 <= r11[2];
cmp204_in1 <= r11[16];
r12[2] <= cmp204_out0;
r12[16] <= cmp204_out1;

cmp205_in0 <= r11[3];
cmp205_in1 <= r11[17];
r12[3] <= cmp205_out0;
r12[17] <= cmp205_out1;

cmp206_in0 <= r11[6];
cmp206_in1 <= r11[20];
r12[6] <= cmp206_out0;
r12[20] <= cmp206_out1;

cmp207_in0 <= r11[7];
cmp207_in1 <= r11[21];
r12[7] <= cmp207_out0;
r12[21] <= cmp207_out1;

cmp208_in0 <= r11[10];
cmp208_in1 <= r11[24];
r12[10] <= cmp208_out0;
r12[24] <= cmp208_out1;

cmp209_in0 <= r11[11];
cmp209_in1 <= r11[25];
r12[11] <= cmp209_out0;
r12[25] <= cmp209_out1;

cmp210_in0 <= r11[14];
cmp210_in1 <= r11[28];
r12[14] <= cmp210_out0;
r12[28] <= cmp210_out1;

cmp211_in0 <= r11[15];
cmp211_in1 <= r11[29];
r12[15] <= cmp211_out0;
r12[29] <= cmp211_out1;

cmp212_in0 <= r11[18];
cmp212_in1 <= r11[32];
r12[18] <= cmp212_out0;
r12[32] <= cmp212_out1;

cmp213_in0 <= r11[19];
cmp213_in1 <= r11[33];
r12[19] <= cmp213_out0;
r12[33] <= cmp213_out1;

cmp214_in0 <= r11[22];
cmp214_in1 <= r11[36];
r12[22] <= cmp214_out0;
r12[36] <= cmp214_out1;

cmp215_in0 <= r11[23];
cmp215_in1 <= r11[37];
r12[23] <= cmp215_out0;
r12[37] <= cmp215_out1;

cmp216_in0 <= r11[26];
cmp216_in1 <= r11[40];
r12[26] <= cmp216_out0;
r12[40] <= cmp216_out1;

cmp217_in0 <= r11[27];
cmp217_in1 <= r11[41];
r12[27] <= cmp217_out0;
r12[41] <= cmp217_out1;

cmp218_in0 <= r11[30];
cmp218_in1 <= r11[44];
r12[30] <= cmp218_out0;
r12[44] <= cmp218_out1;

cmp219_in0 <= r11[31];
cmp219_in1 <= r11[45];
r12[31] <= cmp219_out0;
r12[45] <= cmp219_out1;

cmp220_in0 <= r11[34];
cmp220_in1 <= r11[48];
r12[34] <= cmp220_out0;
r12[48] <= cmp220_out1;

r_12_0_tmp <= r11[0];
r12[0] <= r_12_0_tmp;

r_12_1_tmp <= r11[1];
r12[1] <= r_12_1_tmp;

r_12_4_tmp <= r11[4];
r12[4] <= r_12_4_tmp;

r_12_5_tmp <= r11[5];
r12[5] <= r_12_5_tmp;

r_12_8_tmp <= r11[8];
r12[8] <= r_12_8_tmp;

r_12_9_tmp <= r11[9];
r12[9] <= r_12_9_tmp;

r_12_12_tmp <= r11[12];
r12[12] <= r_12_12_tmp;

r_12_13_tmp <= r11[13];
r12[13] <= r_12_13_tmp;

r_12_35_tmp <= r11[35];
r12[35] <= r_12_35_tmp;

r_12_38_tmp <= r11[38];
r12[38] <= r_12_38_tmp;

r_12_39_tmp <= r11[39];
r12[39] <= r_12_39_tmp;

r_12_42_tmp <= r11[42];
r12[42] <= r_12_42_tmp;

r_12_43_tmp <= r11[43];
r12[43] <= r_12_43_tmp;

r_12_46_tmp <= r11[46];
r12[46] <= r_12_46_tmp;

r_12_47_tmp <= r11[47];
r12[47] <= r_12_47_tmp;

//--------------------------
//---------layer : 13------------
cmp221_in0 <= r12[2];
cmp221_in1 <= r12[8];
r13[2] <= cmp221_out0;
r13[8] <= cmp221_out1;

cmp222_in0 <= r12[3];
cmp222_in1 <= r12[9];
r13[3] <= cmp222_out0;
r13[9] <= cmp222_out1;

cmp223_in0 <= r12[6];
cmp223_in1 <= r12[12];
r13[6] <= cmp223_out0;
r13[12] <= cmp223_out1;

cmp224_in0 <= r12[7];
cmp224_in1 <= r12[13];
r13[7] <= cmp224_out0;
r13[13] <= cmp224_out1;

cmp225_in0 <= r12[10];
cmp225_in1 <= r12[16];
r13[10] <= cmp225_out0;
r13[16] <= cmp225_out1;

cmp226_in0 <= r12[11];
cmp226_in1 <= r12[17];
r13[11] <= cmp226_out0;
r13[17] <= cmp226_out1;

cmp227_in0 <= r12[14];
cmp227_in1 <= r12[20];
r13[14] <= cmp227_out0;
r13[20] <= cmp227_out1;

cmp228_in0 <= r12[15];
cmp228_in1 <= r12[21];
r13[15] <= cmp228_out0;
r13[21] <= cmp228_out1;

cmp229_in0 <= r12[18];
cmp229_in1 <= r12[24];
r13[18] <= cmp229_out0;
r13[24] <= cmp229_out1;

cmp230_in0 <= r12[19];
cmp230_in1 <= r12[25];
r13[19] <= cmp230_out0;
r13[25] <= cmp230_out1;

cmp231_in0 <= r12[22];
cmp231_in1 <= r12[28];
r13[22] <= cmp231_out0;
r13[28] <= cmp231_out1;

cmp232_in0 <= r12[23];
cmp232_in1 <= r12[29];
r13[23] <= cmp232_out0;
r13[29] <= cmp232_out1;

cmp233_in0 <= r12[26];
cmp233_in1 <= r12[32];
r13[26] <= cmp233_out0;
r13[32] <= cmp233_out1;

cmp234_in0 <= r12[27];
cmp234_in1 <= r12[33];
r13[27] <= cmp234_out0;
r13[33] <= cmp234_out1;

cmp235_in0 <= r12[30];
cmp235_in1 <= r12[36];
r13[30] <= cmp235_out0;
r13[36] <= cmp235_out1;

cmp236_in0 <= r12[31];
cmp236_in1 <= r12[37];
r13[31] <= cmp236_out0;
r13[37] <= cmp236_out1;

cmp237_in0 <= r12[34];
cmp237_in1 <= r12[40];
r13[34] <= cmp237_out0;
r13[40] <= cmp237_out1;

cmp238_in0 <= r12[35];
cmp238_in1 <= r12[41];
r13[35] <= cmp238_out0;
r13[41] <= cmp238_out1;

cmp239_in0 <= r12[38];
cmp239_in1 <= r12[44];
r13[38] <= cmp239_out0;
r13[44] <= cmp239_out1;

cmp240_in0 <= r12[39];
cmp240_in1 <= r12[45];
r13[39] <= cmp240_out0;
r13[45] <= cmp240_out1;

cmp241_in0 <= r12[42];
cmp241_in1 <= r12[48];
r13[42] <= cmp241_out0;
r13[48] <= cmp241_out1;

r_13_0_tmp <= r12[0];
r13[0] <= r_13_0_tmp;

r_13_1_tmp <= r12[1];
r13[1] <= r_13_1_tmp;

r_13_4_tmp <= r12[4];
r13[4] <= r_13_4_tmp;

r_13_5_tmp <= r12[5];
r13[5] <= r_13_5_tmp;

r_13_43_tmp <= r12[43];
r13[43] <= r_13_43_tmp;

r_13_46_tmp <= r12[46];
r13[46] <= r_13_46_tmp;

r_13_47_tmp <= r12[47];
r13[47] <= r_13_47_tmp;

//--------------------------
//---------layer : 14------------
cmp242_in0 <= r13[2];
cmp242_in1 <= r13[4];
r14[2] <= cmp242_out0;
r14[4] <= cmp242_out1;

cmp243_in0 <= r13[3];
cmp243_in1 <= r13[5];
r14[3] <= cmp243_out0;
r14[5] <= cmp243_out1;

cmp244_in0 <= r13[6];
cmp244_in1 <= r13[8];
r14[6] <= cmp244_out0;
r14[8] <= cmp244_out1;

cmp245_in0 <= r13[7];
cmp245_in1 <= r13[9];
r14[7] <= cmp245_out0;
r14[9] <= cmp245_out1;

cmp246_in0 <= r13[10];
cmp246_in1 <= r13[12];
r14[10] <= cmp246_out0;
r14[12] <= cmp246_out1;

cmp247_in0 <= r13[11];
cmp247_in1 <= r13[13];
r14[11] <= cmp247_out0;
r14[13] <= cmp247_out1;

cmp248_in0 <= r13[14];
cmp248_in1 <= r13[16];
r14[14] <= cmp248_out0;
r14[16] <= cmp248_out1;

cmp249_in0 <= r13[15];
cmp249_in1 <= r13[17];
r14[15] <= cmp249_out0;
r14[17] <= cmp249_out1;

cmp250_in0 <= r13[18];
cmp250_in1 <= r13[20];
r14[18] <= cmp250_out0;
r14[20] <= cmp250_out1;

cmp251_in0 <= r13[19];
cmp251_in1 <= r13[21];
r14[19] <= cmp251_out0;
r14[21] <= cmp251_out1;

cmp252_in0 <= r13[22];
cmp252_in1 <= r13[24];
r14[22] <= cmp252_out0;
r14[24] <= cmp252_out1;

cmp253_in0 <= r13[23];
cmp253_in1 <= r13[25];
r14[23] <= cmp253_out0;
r14[25] <= cmp253_out1;

cmp254_in0 <= r13[26];
cmp254_in1 <= r13[28];
r14[26] <= cmp254_out0;
r14[28] <= cmp254_out1;

cmp255_in0 <= r13[27];
cmp255_in1 <= r13[29];
r14[27] <= cmp255_out0;
r14[29] <= cmp255_out1;

cmp256_in0 <= r13[30];
cmp256_in1 <= r13[32];
r14[30] <= cmp256_out0;
r14[32] <= cmp256_out1;

cmp257_in0 <= r13[31];
cmp257_in1 <= r13[33];
r14[31] <= cmp257_out0;
r14[33] <= cmp257_out1;

cmp258_in0 <= r13[34];
cmp258_in1 <= r13[36];
r14[34] <= cmp258_out0;
r14[36] <= cmp258_out1;

cmp259_in0 <= r13[35];
cmp259_in1 <= r13[37];
r14[35] <= cmp259_out0;
r14[37] <= cmp259_out1;

cmp260_in0 <= r13[38];
cmp260_in1 <= r13[40];
r14[38] <= cmp260_out0;
r14[40] <= cmp260_out1;

cmp261_in0 <= r13[39];
cmp261_in1 <= r13[41];
r14[39] <= cmp261_out0;
r14[41] <= cmp261_out1;

cmp262_in0 <= r13[42];
cmp262_in1 <= r13[44];
r14[42] <= cmp262_out0;
r14[44] <= cmp262_out1;

cmp263_in0 <= r13[43];
cmp263_in1 <= r13[45];
r14[43] <= cmp263_out0;
r14[45] <= cmp263_out1;

cmp264_in0 <= r13[46];
cmp264_in1 <= r13[48];
r14[46] <= cmp264_out0;
r14[48] <= cmp264_out1;

cmp265_in0 <= r13[0];
cmp265_in1 <= r13[1];
r14[0] <= cmp265_out0;
r14[1] <= cmp265_out1;

r_14_47_tmp <= r13[47];
r14[47] <= r_14_47_tmp;

//--------------------------
//---------layer : 15------------
cmp266_in0 <= r14[2];
cmp266_in1 <= r14[3];
r15[2] <= cmp266_out0;
r15[3] <= cmp266_out1;

cmp267_in0 <= r14[4];
cmp267_in1 <= r14[5];
r15[4] <= cmp267_out0;
r15[5] <= cmp267_out1;

cmp268_in0 <= r14[6];
cmp268_in1 <= r14[7];
r15[6] <= cmp268_out0;
r15[7] <= cmp268_out1;

cmp269_in0 <= r14[8];
cmp269_in1 <= r14[9];
r15[8] <= cmp269_out0;
r15[9] <= cmp269_out1;

cmp270_in0 <= r14[10];
cmp270_in1 <= r14[11];
r15[10] <= cmp270_out0;
r15[11] <= cmp270_out1;

cmp271_in0 <= r14[12];
cmp271_in1 <= r14[13];
r15[12] <= cmp271_out0;
r15[13] <= cmp271_out1;

cmp272_in0 <= r14[14];
cmp272_in1 <= r14[15];
r15[14] <= cmp272_out0;
r15[15] <= cmp272_out1;

cmp273_in0 <= r14[16];
cmp273_in1 <= r14[17];
r15[16] <= cmp273_out0;
r15[17] <= cmp273_out1;

cmp274_in0 <= r14[18];
cmp274_in1 <= r14[19];
r15[18] <= cmp274_out0;
r15[19] <= cmp274_out1;

cmp275_in0 <= r14[20];
cmp275_in1 <= r14[21];
r15[20] <= cmp275_out0;
r15[21] <= cmp275_out1;

cmp276_in0 <= r14[22];
cmp276_in1 <= r14[23];
r15[22] <= cmp276_out0;
r15[23] <= cmp276_out1;

cmp277_in0 <= r14[24];
cmp277_in1 <= r14[25];
r15[24] <= cmp277_out0;
r15[25] <= cmp277_out1;

cmp278_in0 <= r14[26];
cmp278_in1 <= r14[27];
r15[26] <= cmp278_out0;
r15[27] <= cmp278_out1;

cmp279_in0 <= r14[28];
cmp279_in1 <= r14[29];
r15[28] <= cmp279_out0;
r15[29] <= cmp279_out1;

cmp280_in0 <= r14[30];
cmp280_in1 <= r14[31];
r15[30] <= cmp280_out0;
r15[31] <= cmp280_out1;

cmp281_in0 <= r14[32];
cmp281_in1 <= r14[33];
r15[32] <= cmp281_out0;
r15[33] <= cmp281_out1;

cmp282_in0 <= r14[34];
cmp282_in1 <= r14[35];
r15[34] <= cmp282_out0;
r15[35] <= cmp282_out1;

cmp283_in0 <= r14[36];
cmp283_in1 <= r14[37];
r15[36] <= cmp283_out0;
r15[37] <= cmp283_out1;

cmp284_in0 <= r14[38];
cmp284_in1 <= r14[39];
r15[38] <= cmp284_out0;
r15[39] <= cmp284_out1;

cmp285_in0 <= r14[40];
cmp285_in1 <= r14[41];
r15[40] <= cmp285_out0;
r15[41] <= cmp285_out1;

cmp286_in0 <= r14[42];
cmp286_in1 <= r14[43];
r15[42] <= cmp286_out0;
r15[43] <= cmp286_out1;

cmp287_in0 <= r14[44];
cmp287_in1 <= r14[45];
r15[44] <= cmp287_out0;
r15[45] <= cmp287_out1;

cmp288_in0 <= r14[46];
cmp288_in1 <= r14[47];
r15[46] <= cmp288_out0;
r15[47] <= cmp288_out1;

r_15_0_tmp <= r14[0];
r15[0] <= r_15_0_tmp;

r_15_1_tmp <= r14[1];
r15[1] <= r_15_1_tmp;

r_15_48_tmp <= r14[48];
r15[48] <= r_15_48_tmp;

//--------------------------
//---------layer : 16------------
cmp289_in0 <= r15[1];
cmp289_in1 <= r15[32];
r16[1] <= cmp289_out0;
r16[32] <= cmp289_out1;

cmp290_in0 <= r15[3];
cmp290_in1 <= r15[34];
r16[3] <= cmp290_out0;
r16[34] <= cmp290_out1;

cmp291_in0 <= r15[5];
cmp291_in1 <= r15[36];
r16[5] <= cmp291_out0;
r16[36] <= cmp291_out1;

cmp292_in0 <= r15[7];
cmp292_in1 <= r15[38];
r16[7] <= cmp292_out0;
r16[38] <= cmp292_out1;

cmp293_in0 <= r15[9];
cmp293_in1 <= r15[40];
r16[9] <= cmp293_out0;
r16[40] <= cmp293_out1;

cmp294_in0 <= r15[11];
cmp294_in1 <= r15[42];
r16[11] <= cmp294_out0;
r16[42] <= cmp294_out1;

cmp295_in0 <= r15[13];
cmp295_in1 <= r15[44];
r16[13] <= cmp295_out0;
r16[44] <= cmp295_out1;

cmp296_in0 <= r15[15];
cmp296_in1 <= r15[46];
r16[15] <= cmp296_out0;
r16[46] <= cmp296_out1;

cmp297_in0 <= r15[17];
cmp297_in1 <= r15[48];
r16[17] <= cmp297_out0;
r16[48] <= cmp297_out1;

r_16_0_tmp <= r15[0];
r16[0] <= r_16_0_tmp;

r_16_2_tmp <= r15[2];
r16[2] <= r_16_2_tmp;

r_16_4_tmp <= r15[4];
r16[4] <= r_16_4_tmp;

r_16_6_tmp <= r15[6];
r16[6] <= r_16_6_tmp;

r_16_8_tmp <= r15[8];
r16[8] <= r_16_8_tmp;

r_16_10_tmp <= r15[10];
r16[10] <= r_16_10_tmp;

r_16_12_tmp <= r15[12];
r16[12] <= r_16_12_tmp;

r_16_14_tmp <= r15[14];
r16[14] <= r_16_14_tmp;

r_16_16_tmp <= r15[16];
r16[16] <= r_16_16_tmp;

r_16_18_tmp <= r15[18];
r16[18] <= r_16_18_tmp;

r_16_19_tmp <= r15[19];
r16[19] <= r_16_19_tmp;

r_16_20_tmp <= r15[20];
r16[20] <= r_16_20_tmp;

r_16_21_tmp <= r15[21];
r16[21] <= r_16_21_tmp;

r_16_22_tmp <= r15[22];
r16[22] <= r_16_22_tmp;

r_16_23_tmp <= r15[23];
r16[23] <= r_16_23_tmp;

r_16_24_tmp <= r15[24];
r16[24] <= r_16_24_tmp;

r_16_25_tmp <= r15[25];
r16[25] <= r_16_25_tmp;

r_16_26_tmp <= r15[26];
r16[26] <= r_16_26_tmp;

r_16_27_tmp <= r15[27];
r16[27] <= r_16_27_tmp;

r_16_28_tmp <= r15[28];
r16[28] <= r_16_28_tmp;

r_16_29_tmp <= r15[29];
r16[29] <= r_16_29_tmp;

r_16_30_tmp <= r15[30];
r16[30] <= r_16_30_tmp;

r_16_31_tmp <= r15[31];
r16[31] <= r_16_31_tmp;

r_16_33_tmp <= r15[33];
r16[33] <= r_16_33_tmp;

r_16_35_tmp <= r15[35];
r16[35] <= r_16_35_tmp;

r_16_37_tmp <= r15[37];
r16[37] <= r_16_37_tmp;

r_16_39_tmp <= r15[39];
r16[39] <= r_16_39_tmp;

r_16_41_tmp <= r15[41];
r16[41] <= r_16_41_tmp;

r_16_43_tmp <= r15[43];
r16[43] <= r_16_43_tmp;

r_16_45_tmp <= r15[45];
r16[45] <= r_16_45_tmp;

r_16_47_tmp <= r15[47];
r16[47] <= r_16_47_tmp;

//--------------------------
//---------layer : 17------------
cmp298_in0 <= r16[9];
cmp298_in1 <= r16[24];
r17[9] <= cmp298_out0;
r17[24] <= cmp298_out1;

cmp299_in0 <= r16[11];
cmp299_in1 <= r16[26];
r17[11] <= cmp299_out0;
r17[26] <= cmp299_out1;

cmp300_in0 <= r16[13];
cmp300_in1 <= r16[28];
r17[13] <= cmp300_out0;
r17[28] <= cmp300_out1;

cmp301_in0 <= r16[15];
cmp301_in1 <= r16[30];
r17[15] <= cmp301_out0;
r17[30] <= cmp301_out1;

cmp302_in0 <= r16[17];
cmp302_in1 <= r16[32];
r17[17] <= cmp302_out0;
r17[32] <= cmp302_out1;

cmp303_in0 <= r16[19];
cmp303_in1 <= r16[34];
r17[19] <= cmp303_out0;
r17[34] <= cmp303_out1;

cmp304_in0 <= r16[21];
cmp304_in1 <= r16[36];
r17[21] <= cmp304_out0;
r17[36] <= cmp304_out1;

cmp305_in0 <= r16[23];
cmp305_in1 <= r16[38];
r17[23] <= cmp305_out0;
r17[38] <= cmp305_out1;

r_17_0_tmp <= r16[0];
r17[0] <= r_17_0_tmp;

r_17_1_tmp <= r16[1];
r17[1] <= r_17_1_tmp;

r_17_2_tmp <= r16[2];
r17[2] <= r_17_2_tmp;

r_17_3_tmp <= r16[3];
r17[3] <= r_17_3_tmp;

r_17_4_tmp <= r16[4];
r17[4] <= r_17_4_tmp;

r_17_5_tmp <= r16[5];
r17[5] <= r_17_5_tmp;

r_17_6_tmp <= r16[6];
r17[6] <= r_17_6_tmp;

r_17_7_tmp <= r16[7];
r17[7] <= r_17_7_tmp;

r_17_8_tmp <= r16[8];
r17[8] <= r_17_8_tmp;

r_17_10_tmp <= r16[10];
r17[10] <= r_17_10_tmp;

r_17_12_tmp <= r16[12];
r17[12] <= r_17_12_tmp;

r_17_14_tmp <= r16[14];
r17[14] <= r_17_14_tmp;

r_17_16_tmp <= r16[16];
r17[16] <= r_17_16_tmp;

r_17_18_tmp <= r16[18];
r17[18] <= r_17_18_tmp;

r_17_20_tmp <= r16[20];
r17[20] <= r_17_20_tmp;

r_17_22_tmp <= r16[22];
r17[22] <= r_17_22_tmp;

r_17_25_tmp <= r16[25];
r17[25] <= r_17_25_tmp;

r_17_27_tmp <= r16[27];
r17[27] <= r_17_27_tmp;

r_17_29_tmp <= r16[29];
r17[29] <= r_17_29_tmp;

r_17_31_tmp <= r16[31];
r17[31] <= r_17_31_tmp;

r_17_33_tmp <= r16[33];
r17[33] <= r_17_33_tmp;

r_17_35_tmp <= r16[35];
r17[35] <= r_17_35_tmp;

r_17_37_tmp <= r16[37];
r17[37] <= r_17_37_tmp;

r_17_39_tmp <= r16[39];
r17[39] <= r_17_39_tmp;

r_17_40_tmp <= r16[40];
r17[40] <= r_17_40_tmp;

r_17_41_tmp <= r16[41];
r17[41] <= r_17_41_tmp;

r_17_42_tmp <= r16[42];
r17[42] <= r_17_42_tmp;

r_17_43_tmp <= r16[43];
r17[43] <= r_17_43_tmp;

r_17_44_tmp <= r16[44];
r17[44] <= r_17_44_tmp;

r_17_45_tmp <= r16[45];
r17[45] <= r_17_45_tmp;

r_17_46_tmp <= r16[46];
r17[46] <= r_17_46_tmp;

r_17_47_tmp <= r16[47];
r17[47] <= r_17_47_tmp;

r_17_48_tmp <= r16[48];
r17[48] <= r_17_48_tmp;

//--------------------------
//---------layer : 18------------
cmp306_in0 <= r17[17];
cmp306_in1 <= r17[24];
r18[17] <= cmp306_out0;
r18[24] <= cmp306_out1;

cmp307_in0 <= r17[19];
cmp307_in1 <= r17[26];
r18[19] <= cmp307_out0;
r18[26] <= cmp307_out1;

cmp308_in0 <= r17[21];
cmp308_in1 <= r17[28];
r18[21] <= cmp308_out0;
r18[28] <= cmp308_out1;

cmp309_in0 <= r17[23];
cmp309_in1 <= r17[30];
r18[23] <= cmp309_out0;
r18[30] <= cmp309_out1;

r_18_0_tmp <= r17[0];
r18[0] <= r_18_0_tmp;

r_18_1_tmp <= r17[1];
r18[1] <= r_18_1_tmp;

r_18_2_tmp <= r17[2];
r18[2] <= r_18_2_tmp;

r_18_3_tmp <= r17[3];
r18[3] <= r_18_3_tmp;

r_18_4_tmp <= r17[4];
r18[4] <= r_18_4_tmp;

r_18_5_tmp <= r17[5];
r18[5] <= r_18_5_tmp;

r_18_6_tmp <= r17[6];
r18[6] <= r_18_6_tmp;

r_18_7_tmp <= r17[7];
r18[7] <= r_18_7_tmp;

r_18_8_tmp <= r17[8];
r18[8] <= r_18_8_tmp;

r_18_9_tmp <= r17[9];
r18[9] <= r_18_9_tmp;

r_18_10_tmp <= r17[10];
r18[10] <= r_18_10_tmp;

r_18_11_tmp <= r17[11];
r18[11] <= r_18_11_tmp;

r_18_12_tmp <= r17[12];
r18[12] <= r_18_12_tmp;

r_18_13_tmp <= r17[13];
r18[13] <= r_18_13_tmp;

r_18_14_tmp <= r17[14];
r18[14] <= r_18_14_tmp;

r_18_15_tmp <= r17[15];
r18[15] <= r_18_15_tmp;

r_18_16_tmp <= r17[16];
r18[16] <= r_18_16_tmp;

r_18_18_tmp <= r17[18];
r18[18] <= r_18_18_tmp;

r_18_20_tmp <= r17[20];
r18[20] <= r_18_20_tmp;

r_18_22_tmp <= r17[22];
r18[22] <= r_18_22_tmp;

r_18_25_tmp <= r17[25];
r18[25] <= r_18_25_tmp;

r_18_27_tmp <= r17[27];
r18[27] <= r_18_27_tmp;

r_18_29_tmp <= r17[29];
r18[29] <= r_18_29_tmp;

r_18_31_tmp <= r17[31];
r18[31] <= r_18_31_tmp;

r_18_32_tmp <= r17[32];
r18[32] <= r_18_32_tmp;

r_18_33_tmp <= r17[33];
r18[33] <= r_18_33_tmp;

r_18_34_tmp <= r17[34];
r18[34] <= r_18_34_tmp;

r_18_35_tmp <= r17[35];
r18[35] <= r_18_35_tmp;

r_18_36_tmp <= r17[36];
r18[36] <= r_18_36_tmp;

r_18_37_tmp <= r17[37];
r18[37] <= r_18_37_tmp;

r_18_38_tmp <= r17[38];
r18[38] <= r_18_38_tmp;

r_18_39_tmp <= r17[39];
r18[39] <= r_18_39_tmp;

r_18_40_tmp <= r17[40];
r18[40] <= r_18_40_tmp;

r_18_41_tmp <= r17[41];
r18[41] <= r_18_41_tmp;

r_18_42_tmp <= r17[42];
r18[42] <= r_18_42_tmp;

r_18_43_tmp <= r17[43];
r18[43] <= r_18_43_tmp;

r_18_44_tmp <= r17[44];
r18[44] <= r_18_44_tmp;

r_18_45_tmp <= r17[45];
r18[45] <= r_18_45_tmp;

r_18_46_tmp <= r17[46];
r18[46] <= r_18_46_tmp;

r_18_47_tmp <= r17[47];
r18[47] <= r_18_47_tmp;

r_18_48_tmp <= r17[48];
r18[48] <= r_18_48_tmp;

//--------------------------
//---------layer : 19------------
cmp310_in0 <= r18[21];
cmp310_in1 <= r18[24];
r19[21] <= cmp310_out0;
r19[24] <= cmp310_out1;

cmp311_in0 <= r18[23];
cmp311_in1 <= r18[26];
r19[23] <= cmp311_out0;
r19[26] <= cmp311_out1;

r_19_0_tmp <= r18[0];
r19[0] <= r_19_0_tmp;

r_19_1_tmp <= r18[1];
r19[1] <= r_19_1_tmp;

r_19_2_tmp <= r18[2];
r19[2] <= r_19_2_tmp;

r_19_3_tmp <= r18[3];
r19[3] <= r_19_3_tmp;

r_19_4_tmp <= r18[4];
r19[4] <= r_19_4_tmp;

r_19_5_tmp <= r18[5];
r19[5] <= r_19_5_tmp;

r_19_6_tmp <= r18[6];
r19[6] <= r_19_6_tmp;

r_19_7_tmp <= r18[7];
r19[7] <= r_19_7_tmp;

r_19_8_tmp <= r18[8];
r19[8] <= r_19_8_tmp;

r_19_9_tmp <= r18[9];
r19[9] <= r_19_9_tmp;

r_19_10_tmp <= r18[10];
r19[10] <= r_19_10_tmp;

r_19_11_tmp <= r18[11];
r19[11] <= r_19_11_tmp;

r_19_12_tmp <= r18[12];
r19[12] <= r_19_12_tmp;

r_19_13_tmp <= r18[13];
r19[13] <= r_19_13_tmp;

r_19_14_tmp <= r18[14];
r19[14] <= r_19_14_tmp;

r_19_15_tmp <= r18[15];
r19[15] <= r_19_15_tmp;

r_19_16_tmp <= r18[16];
r19[16] <= r_19_16_tmp;

r_19_17_tmp <= r18[17];
r19[17] <= r_19_17_tmp;

r_19_18_tmp <= r18[18];
r19[18] <= r_19_18_tmp;

r_19_19_tmp <= r18[19];
r19[19] <= r_19_19_tmp;

r_19_20_tmp <= r18[20];
r19[20] <= r_19_20_tmp;

r_19_22_tmp <= r18[22];
r19[22] <= r_19_22_tmp;

r_19_25_tmp <= r18[25];
r19[25] <= r_19_25_tmp;

r_19_27_tmp <= r18[27];
r19[27] <= r_19_27_tmp;

r_19_28_tmp <= r18[28];
r19[28] <= r_19_28_tmp;

r_19_29_tmp <= r18[29];
r19[29] <= r_19_29_tmp;

r_19_30_tmp <= r18[30];
r19[30] <= r_19_30_tmp;

r_19_31_tmp <= r18[31];
r19[31] <= r_19_31_tmp;

r_19_32_tmp <= r18[32];
r19[32] <= r_19_32_tmp;

r_19_33_tmp <= r18[33];
r19[33] <= r_19_33_tmp;

r_19_34_tmp <= r18[34];
r19[34] <= r_19_34_tmp;

r_19_35_tmp <= r18[35];
r19[35] <= r_19_35_tmp;

r_19_36_tmp <= r18[36];
r19[36] <= r_19_36_tmp;

r_19_37_tmp <= r18[37];
r19[37] <= r_19_37_tmp;

r_19_38_tmp <= r18[38];
r19[38] <= r_19_38_tmp;

r_19_39_tmp <= r18[39];
r19[39] <= r_19_39_tmp;

r_19_40_tmp <= r18[40];
r19[40] <= r_19_40_tmp;

r_19_41_tmp <= r18[41];
r19[41] <= r_19_41_tmp;

r_19_42_tmp <= r18[42];
r19[42] <= r_19_42_tmp;

r_19_43_tmp <= r18[43];
r19[43] <= r_19_43_tmp;

r_19_44_tmp <= r18[44];
r19[44] <= r_19_44_tmp;

r_19_45_tmp <= r18[45];
r19[45] <= r_19_45_tmp;

r_19_46_tmp <= r18[46];
r19[46] <= r_19_46_tmp;

r_19_47_tmp <= r18[47];
r19[47] <= r_19_47_tmp;

r_19_48_tmp <= r18[48];
r19[48] <= r_19_48_tmp;

//--------------------------
//---------layer : 20------------
cmp312_in0 <= r19[23];
cmp312_in1 <= r19[24];
r20[23] <= cmp312_out0;
r20[24] <= cmp312_out1;

r_20_0_tmp <= r19[0];
r20[0] <= r_20_0_tmp;

r_20_1_tmp <= r19[1];
r20[1] <= r_20_1_tmp;

r_20_2_tmp <= r19[2];
r20[2] <= r_20_2_tmp;

r_20_3_tmp <= r19[3];
r20[3] <= r_20_3_tmp;

r_20_4_tmp <= r19[4];
r20[4] <= r_20_4_tmp;

r_20_5_tmp <= r19[5];
r20[5] <= r_20_5_tmp;

r_20_6_tmp <= r19[6];
r20[6] <= r_20_6_tmp;

r_20_7_tmp <= r19[7];
r20[7] <= r_20_7_tmp;

r_20_8_tmp <= r19[8];
r20[8] <= r_20_8_tmp;

r_20_9_tmp <= r19[9];
r20[9] <= r_20_9_tmp;

r_20_10_tmp <= r19[10];
r20[10] <= r_20_10_tmp;

r_20_11_tmp <= r19[11];
r20[11] <= r_20_11_tmp;

r_20_12_tmp <= r19[12];
r20[12] <= r_20_12_tmp;

r_20_13_tmp <= r19[13];
r20[13] <= r_20_13_tmp;

r_20_14_tmp <= r19[14];
r20[14] <= r_20_14_tmp;

r_20_15_tmp <= r19[15];
r20[15] <= r_20_15_tmp;

r_20_16_tmp <= r19[16];
r20[16] <= r_20_16_tmp;

r_20_17_tmp <= r19[17];
r20[17] <= r_20_17_tmp;

r_20_18_tmp <= r19[18];
r20[18] <= r_20_18_tmp;

r_20_19_tmp <= r19[19];
r20[19] <= r_20_19_tmp;

r_20_20_tmp <= r19[20];
r20[20] <= r_20_20_tmp;

r_20_21_tmp <= r19[21];
r20[21] <= r_20_21_tmp;

r_20_22_tmp <= r19[22];
r20[22] <= r_20_22_tmp;

r_20_25_tmp <= r19[25];
r20[25] <= r_20_25_tmp;

r_20_26_tmp <= r19[26];
r20[26] <= r_20_26_tmp;

r_20_27_tmp <= r19[27];
r20[27] <= r_20_27_tmp;

r_20_28_tmp <= r19[28];
r20[28] <= r_20_28_tmp;

r_20_29_tmp <= r19[29];
r20[29] <= r_20_29_tmp;

r_20_30_tmp <= r19[30];
r20[30] <= r_20_30_tmp;

r_20_31_tmp <= r19[31];
r20[31] <= r_20_31_tmp;

r_20_32_tmp <= r19[32];
r20[32] <= r_20_32_tmp;

r_20_33_tmp <= r19[33];
r20[33] <= r_20_33_tmp;

r_20_34_tmp <= r19[34];
r20[34] <= r_20_34_tmp;

r_20_35_tmp <= r19[35];
r20[35] <= r_20_35_tmp;

r_20_36_tmp <= r19[36];
r20[36] <= r_20_36_tmp;

r_20_37_tmp <= r19[37];
r20[37] <= r_20_37_tmp;

r_20_38_tmp <= r19[38];
r20[38] <= r_20_38_tmp;

r_20_39_tmp <= r19[39];
r20[39] <= r_20_39_tmp;

r_20_40_tmp <= r19[40];
r20[40] <= r_20_40_tmp;

r_20_41_tmp <= r19[41];
r20[41] <= r_20_41_tmp;

r_20_42_tmp <= r19[42];
r20[42] <= r_20_42_tmp;

r_20_43_tmp <= r19[43];
r20[43] <= r_20_43_tmp;

r_20_44_tmp <= r19[44];
r20[44] <= r_20_44_tmp;

r_20_45_tmp <= r19[45];
r20[45] <= r_20_45_tmp;

r_20_46_tmp <= r19[46];
r20[46] <= r_20_46_tmp;

r_20_47_tmp <= r19[47];
r20[47] <= r_20_47_tmp;

r_20_48_tmp <= r19[48];
r20[48] <= r_20_48_tmp;

//--------------------------
end
cmp cmp0 (.in0(cmp0_in0), .in1(cmp0_in1), .out0(cmp0_out0), .out1(cmp0_out1));
cmp cmp1 (.in0(cmp1_in0), .in1(cmp1_in1), .out0(cmp1_out0), .out1(cmp1_out1));
cmp cmp2 (.in0(cmp2_in0), .in1(cmp2_in1), .out0(cmp2_out0), .out1(cmp2_out1));
cmp cmp3 (.in0(cmp3_in0), .in1(cmp3_in1), .out0(cmp3_out0), .out1(cmp3_out1));
cmp cmp4 (.in0(cmp4_in0), .in1(cmp4_in1), .out0(cmp4_out0), .out1(cmp4_out1));
cmp cmp5 (.in0(cmp5_in0), .in1(cmp5_in1), .out0(cmp5_out0), .out1(cmp5_out1));
cmp cmp6 (.in0(cmp6_in0), .in1(cmp6_in1), .out0(cmp6_out0), .out1(cmp6_out1));
cmp cmp7 (.in0(cmp7_in0), .in1(cmp7_in1), .out0(cmp7_out0), .out1(cmp7_out1));
cmp cmp8 (.in0(cmp8_in0), .in1(cmp8_in1), .out0(cmp8_out0), .out1(cmp8_out1));
cmp cmp9 (.in0(cmp9_in0), .in1(cmp9_in1), .out0(cmp9_out0), .out1(cmp9_out1));
cmp cmp10 (.in0(cmp10_in0), .in1(cmp10_in1), .out0(cmp10_out0), .out1(cmp10_out1));
cmp cmp11 (.in0(cmp11_in0), .in1(cmp11_in1), .out0(cmp11_out0), .out1(cmp11_out1));
cmp cmp12 (.in0(cmp12_in0), .in1(cmp12_in1), .out0(cmp12_out0), .out1(cmp12_out1));
cmp cmp13 (.in0(cmp13_in0), .in1(cmp13_in1), .out0(cmp13_out0), .out1(cmp13_out1));
cmp cmp14 (.in0(cmp14_in0), .in1(cmp14_in1), .out0(cmp14_out0), .out1(cmp14_out1));
cmp cmp15 (.in0(cmp15_in0), .in1(cmp15_in1), .out0(cmp15_out0), .out1(cmp15_out1));
cmp cmp16 (.in0(cmp16_in0), .in1(cmp16_in1), .out0(cmp16_out0), .out1(cmp16_out1));
cmp cmp17 (.in0(cmp17_in0), .in1(cmp17_in1), .out0(cmp17_out0), .out1(cmp17_out1));
cmp cmp18 (.in0(cmp18_in0), .in1(cmp18_in1), .out0(cmp18_out0), .out1(cmp18_out1));
cmp cmp19 (.in0(cmp19_in0), .in1(cmp19_in1), .out0(cmp19_out0), .out1(cmp19_out1));
cmp cmp20 (.in0(cmp20_in0), .in1(cmp20_in1), .out0(cmp20_out0), .out1(cmp20_out1));
cmp cmp21 (.in0(cmp21_in0), .in1(cmp21_in1), .out0(cmp21_out0), .out1(cmp21_out1));
cmp cmp22 (.in0(cmp22_in0), .in1(cmp22_in1), .out0(cmp22_out0), .out1(cmp22_out1));
cmp cmp23 (.in0(cmp23_in0), .in1(cmp23_in1), .out0(cmp23_out0), .out1(cmp23_out1));
cmp cmp24 (.in0(cmp24_in0), .in1(cmp24_in1), .out0(cmp24_out0), .out1(cmp24_out1));
cmp cmp25 (.in0(cmp25_in0), .in1(cmp25_in1), .out0(cmp25_out0), .out1(cmp25_out1));
cmp cmp26 (.in0(cmp26_in0), .in1(cmp26_in1), .out0(cmp26_out0), .out1(cmp26_out1));
cmp cmp27 (.in0(cmp27_in0), .in1(cmp27_in1), .out0(cmp27_out0), .out1(cmp27_out1));
cmp cmp28 (.in0(cmp28_in0), .in1(cmp28_in1), .out0(cmp28_out0), .out1(cmp28_out1));
cmp cmp29 (.in0(cmp29_in0), .in1(cmp29_in1), .out0(cmp29_out0), .out1(cmp29_out1));
cmp cmp30 (.in0(cmp30_in0), .in1(cmp30_in1), .out0(cmp30_out0), .out1(cmp30_out1));
cmp cmp31 (.in0(cmp31_in0), .in1(cmp31_in1), .out0(cmp31_out0), .out1(cmp31_out1));
cmp cmp32 (.in0(cmp32_in0), .in1(cmp32_in1), .out0(cmp32_out0), .out1(cmp32_out1));
cmp cmp33 (.in0(cmp33_in0), .in1(cmp33_in1), .out0(cmp33_out0), .out1(cmp33_out1));
cmp cmp34 (.in0(cmp34_in0), .in1(cmp34_in1), .out0(cmp34_out0), .out1(cmp34_out1));
cmp cmp35 (.in0(cmp35_in0), .in1(cmp35_in1), .out0(cmp35_out0), .out1(cmp35_out1));
cmp cmp36 (.in0(cmp36_in0), .in1(cmp36_in1), .out0(cmp36_out0), .out1(cmp36_out1));
cmp cmp37 (.in0(cmp37_in0), .in1(cmp37_in1), .out0(cmp37_out0), .out1(cmp37_out1));
cmp cmp38 (.in0(cmp38_in0), .in1(cmp38_in1), .out0(cmp38_out0), .out1(cmp38_out1));
cmp cmp39 (.in0(cmp39_in0), .in1(cmp39_in1), .out0(cmp39_out0), .out1(cmp39_out1));
cmp cmp40 (.in0(cmp40_in0), .in1(cmp40_in1), .out0(cmp40_out0), .out1(cmp40_out1));
cmp cmp41 (.in0(cmp41_in0), .in1(cmp41_in1), .out0(cmp41_out0), .out1(cmp41_out1));
cmp cmp42 (.in0(cmp42_in0), .in1(cmp42_in1), .out0(cmp42_out0), .out1(cmp42_out1));
cmp cmp43 (.in0(cmp43_in0), .in1(cmp43_in1), .out0(cmp43_out0), .out1(cmp43_out1));
cmp cmp44 (.in0(cmp44_in0), .in1(cmp44_in1), .out0(cmp44_out0), .out1(cmp44_out1));
cmp cmp45 (.in0(cmp45_in0), .in1(cmp45_in1), .out0(cmp45_out0), .out1(cmp45_out1));
cmp cmp46 (.in0(cmp46_in0), .in1(cmp46_in1), .out0(cmp46_out0), .out1(cmp46_out1));
cmp cmp47 (.in0(cmp47_in0), .in1(cmp47_in1), .out0(cmp47_out0), .out1(cmp47_out1));
cmp cmp48 (.in0(cmp48_in0), .in1(cmp48_in1), .out0(cmp48_out0), .out1(cmp48_out1));
cmp cmp49 (.in0(cmp49_in0), .in1(cmp49_in1), .out0(cmp49_out0), .out1(cmp49_out1));
cmp cmp50 (.in0(cmp50_in0), .in1(cmp50_in1), .out0(cmp50_out0), .out1(cmp50_out1));
cmp cmp51 (.in0(cmp51_in0), .in1(cmp51_in1), .out0(cmp51_out0), .out1(cmp51_out1));
cmp cmp52 (.in0(cmp52_in0), .in1(cmp52_in1), .out0(cmp52_out0), .out1(cmp52_out1));
cmp cmp53 (.in0(cmp53_in0), .in1(cmp53_in1), .out0(cmp53_out0), .out1(cmp53_out1));
cmp cmp54 (.in0(cmp54_in0), .in1(cmp54_in1), .out0(cmp54_out0), .out1(cmp54_out1));
cmp cmp55 (.in0(cmp55_in0), .in1(cmp55_in1), .out0(cmp55_out0), .out1(cmp55_out1));
cmp cmp56 (.in0(cmp56_in0), .in1(cmp56_in1), .out0(cmp56_out0), .out1(cmp56_out1));
cmp cmp57 (.in0(cmp57_in0), .in1(cmp57_in1), .out0(cmp57_out0), .out1(cmp57_out1));
cmp cmp58 (.in0(cmp58_in0), .in1(cmp58_in1), .out0(cmp58_out0), .out1(cmp58_out1));
cmp cmp59 (.in0(cmp59_in0), .in1(cmp59_in1), .out0(cmp59_out0), .out1(cmp59_out1));
cmp cmp60 (.in0(cmp60_in0), .in1(cmp60_in1), .out0(cmp60_out0), .out1(cmp60_out1));
cmp cmp61 (.in0(cmp61_in0), .in1(cmp61_in1), .out0(cmp61_out0), .out1(cmp61_out1));
cmp cmp62 (.in0(cmp62_in0), .in1(cmp62_in1), .out0(cmp62_out0), .out1(cmp62_out1));
cmp cmp63 (.in0(cmp63_in0), .in1(cmp63_in1), .out0(cmp63_out0), .out1(cmp63_out1));
cmp cmp64 (.in0(cmp64_in0), .in1(cmp64_in1), .out0(cmp64_out0), .out1(cmp64_out1));
cmp cmp65 (.in0(cmp65_in0), .in1(cmp65_in1), .out0(cmp65_out0), .out1(cmp65_out1));
cmp cmp66 (.in0(cmp66_in0), .in1(cmp66_in1), .out0(cmp66_out0), .out1(cmp66_out1));
cmp cmp67 (.in0(cmp67_in0), .in1(cmp67_in1), .out0(cmp67_out0), .out1(cmp67_out1));
cmp cmp68 (.in0(cmp68_in0), .in1(cmp68_in1), .out0(cmp68_out0), .out1(cmp68_out1));
cmp cmp69 (.in0(cmp69_in0), .in1(cmp69_in1), .out0(cmp69_out0), .out1(cmp69_out1));
cmp cmp70 (.in0(cmp70_in0), .in1(cmp70_in1), .out0(cmp70_out0), .out1(cmp70_out1));
cmp cmp71 (.in0(cmp71_in0), .in1(cmp71_in1), .out0(cmp71_out0), .out1(cmp71_out1));
cmp cmp72 (.in0(cmp72_in0), .in1(cmp72_in1), .out0(cmp72_out0), .out1(cmp72_out1));
cmp cmp73 (.in0(cmp73_in0), .in1(cmp73_in1), .out0(cmp73_out0), .out1(cmp73_out1));
cmp cmp74 (.in0(cmp74_in0), .in1(cmp74_in1), .out0(cmp74_out0), .out1(cmp74_out1));
cmp cmp75 (.in0(cmp75_in0), .in1(cmp75_in1), .out0(cmp75_out0), .out1(cmp75_out1));
cmp cmp76 (.in0(cmp76_in0), .in1(cmp76_in1), .out0(cmp76_out0), .out1(cmp76_out1));
cmp cmp77 (.in0(cmp77_in0), .in1(cmp77_in1), .out0(cmp77_out0), .out1(cmp77_out1));
cmp cmp78 (.in0(cmp78_in0), .in1(cmp78_in1), .out0(cmp78_out0), .out1(cmp78_out1));
cmp cmp79 (.in0(cmp79_in0), .in1(cmp79_in1), .out0(cmp79_out0), .out1(cmp79_out1));
cmp cmp80 (.in0(cmp80_in0), .in1(cmp80_in1), .out0(cmp80_out0), .out1(cmp80_out1));
cmp cmp81 (.in0(cmp81_in0), .in1(cmp81_in1), .out0(cmp81_out0), .out1(cmp81_out1));
cmp cmp82 (.in0(cmp82_in0), .in1(cmp82_in1), .out0(cmp82_out0), .out1(cmp82_out1));
cmp cmp83 (.in0(cmp83_in0), .in1(cmp83_in1), .out0(cmp83_out0), .out1(cmp83_out1));
cmp cmp84 (.in0(cmp84_in0), .in1(cmp84_in1), .out0(cmp84_out0), .out1(cmp84_out1));
cmp cmp85 (.in0(cmp85_in0), .in1(cmp85_in1), .out0(cmp85_out0), .out1(cmp85_out1));
cmp cmp86 (.in0(cmp86_in0), .in1(cmp86_in1), .out0(cmp86_out0), .out1(cmp86_out1));
cmp cmp87 (.in0(cmp87_in0), .in1(cmp87_in1), .out0(cmp87_out0), .out1(cmp87_out1));
cmp cmp88 (.in0(cmp88_in0), .in1(cmp88_in1), .out0(cmp88_out0), .out1(cmp88_out1));
cmp cmp89 (.in0(cmp89_in0), .in1(cmp89_in1), .out0(cmp89_out0), .out1(cmp89_out1));
cmp cmp90 (.in0(cmp90_in0), .in1(cmp90_in1), .out0(cmp90_out0), .out1(cmp90_out1));
cmp cmp91 (.in0(cmp91_in0), .in1(cmp91_in1), .out0(cmp91_out0), .out1(cmp91_out1));
cmp cmp92 (.in0(cmp92_in0), .in1(cmp92_in1), .out0(cmp92_out0), .out1(cmp92_out1));
cmp cmp93 (.in0(cmp93_in0), .in1(cmp93_in1), .out0(cmp93_out0), .out1(cmp93_out1));
cmp cmp94 (.in0(cmp94_in0), .in1(cmp94_in1), .out0(cmp94_out0), .out1(cmp94_out1));
cmp cmp95 (.in0(cmp95_in0), .in1(cmp95_in1), .out0(cmp95_out0), .out1(cmp95_out1));
cmp cmp96 (.in0(cmp96_in0), .in1(cmp96_in1), .out0(cmp96_out0), .out1(cmp96_out1));
cmp cmp97 (.in0(cmp97_in0), .in1(cmp97_in1), .out0(cmp97_out0), .out1(cmp97_out1));
cmp cmp98 (.in0(cmp98_in0), .in1(cmp98_in1), .out0(cmp98_out0), .out1(cmp98_out1));
cmp cmp99 (.in0(cmp99_in0), .in1(cmp99_in1), .out0(cmp99_out0), .out1(cmp99_out1));
cmp cmp100 (.in0(cmp100_in0), .in1(cmp100_in1), .out0(cmp100_out0), .out1(cmp100_out1));
cmp cmp101 (.in0(cmp101_in0), .in1(cmp101_in1), .out0(cmp101_out0), .out1(cmp101_out1));
cmp cmp102 (.in0(cmp102_in0), .in1(cmp102_in1), .out0(cmp102_out0), .out1(cmp102_out1));
cmp cmp103 (.in0(cmp103_in0), .in1(cmp103_in1), .out0(cmp103_out0), .out1(cmp103_out1));
cmp cmp104 (.in0(cmp104_in0), .in1(cmp104_in1), .out0(cmp104_out0), .out1(cmp104_out1));
cmp cmp105 (.in0(cmp105_in0), .in1(cmp105_in1), .out0(cmp105_out0), .out1(cmp105_out1));
cmp cmp106 (.in0(cmp106_in0), .in1(cmp106_in1), .out0(cmp106_out0), .out1(cmp106_out1));
cmp cmp107 (.in0(cmp107_in0), .in1(cmp107_in1), .out0(cmp107_out0), .out1(cmp107_out1));
cmp cmp108 (.in0(cmp108_in0), .in1(cmp108_in1), .out0(cmp108_out0), .out1(cmp108_out1));
cmp cmp109 (.in0(cmp109_in0), .in1(cmp109_in1), .out0(cmp109_out0), .out1(cmp109_out1));
cmp cmp110 (.in0(cmp110_in0), .in1(cmp110_in1), .out0(cmp110_out0), .out1(cmp110_out1));
cmp cmp111 (.in0(cmp111_in0), .in1(cmp111_in1), .out0(cmp111_out0), .out1(cmp111_out1));
cmp cmp112 (.in0(cmp112_in0), .in1(cmp112_in1), .out0(cmp112_out0), .out1(cmp112_out1));
cmp cmp113 (.in0(cmp113_in0), .in1(cmp113_in1), .out0(cmp113_out0), .out1(cmp113_out1));
cmp cmp114 (.in0(cmp114_in0), .in1(cmp114_in1), .out0(cmp114_out0), .out1(cmp114_out1));
cmp cmp115 (.in0(cmp115_in0), .in1(cmp115_in1), .out0(cmp115_out0), .out1(cmp115_out1));
cmp cmp116 (.in0(cmp116_in0), .in1(cmp116_in1), .out0(cmp116_out0), .out1(cmp116_out1));
cmp cmp117 (.in0(cmp117_in0), .in1(cmp117_in1), .out0(cmp117_out0), .out1(cmp117_out1));
cmp cmp118 (.in0(cmp118_in0), .in1(cmp118_in1), .out0(cmp118_out0), .out1(cmp118_out1));
cmp cmp119 (.in0(cmp119_in0), .in1(cmp119_in1), .out0(cmp119_out0), .out1(cmp119_out1));
cmp cmp120 (.in0(cmp120_in0), .in1(cmp120_in1), .out0(cmp120_out0), .out1(cmp120_out1));
cmp cmp121 (.in0(cmp121_in0), .in1(cmp121_in1), .out0(cmp121_out0), .out1(cmp121_out1));
cmp cmp122 (.in0(cmp122_in0), .in1(cmp122_in1), .out0(cmp122_out0), .out1(cmp122_out1));
cmp cmp123 (.in0(cmp123_in0), .in1(cmp123_in1), .out0(cmp123_out0), .out1(cmp123_out1));
cmp cmp124 (.in0(cmp124_in0), .in1(cmp124_in1), .out0(cmp124_out0), .out1(cmp124_out1));
cmp cmp125 (.in0(cmp125_in0), .in1(cmp125_in1), .out0(cmp125_out0), .out1(cmp125_out1));
cmp cmp126 (.in0(cmp126_in0), .in1(cmp126_in1), .out0(cmp126_out0), .out1(cmp126_out1));
cmp cmp127 (.in0(cmp127_in0), .in1(cmp127_in1), .out0(cmp127_out0), .out1(cmp127_out1));
cmp cmp128 (.in0(cmp128_in0), .in1(cmp128_in1), .out0(cmp128_out0), .out1(cmp128_out1));
cmp cmp129 (.in0(cmp129_in0), .in1(cmp129_in1), .out0(cmp129_out0), .out1(cmp129_out1));
cmp cmp130 (.in0(cmp130_in0), .in1(cmp130_in1), .out0(cmp130_out0), .out1(cmp130_out1));
cmp cmp131 (.in0(cmp131_in0), .in1(cmp131_in1), .out0(cmp131_out0), .out1(cmp131_out1));
cmp cmp132 (.in0(cmp132_in0), .in1(cmp132_in1), .out0(cmp132_out0), .out1(cmp132_out1));
cmp cmp133 (.in0(cmp133_in0), .in1(cmp133_in1), .out0(cmp133_out0), .out1(cmp133_out1));
cmp cmp134 (.in0(cmp134_in0), .in1(cmp134_in1), .out0(cmp134_out0), .out1(cmp134_out1));
cmp cmp135 (.in0(cmp135_in0), .in1(cmp135_in1), .out0(cmp135_out0), .out1(cmp135_out1));
cmp cmp136 (.in0(cmp136_in0), .in1(cmp136_in1), .out0(cmp136_out0), .out1(cmp136_out1));
cmp cmp137 (.in0(cmp137_in0), .in1(cmp137_in1), .out0(cmp137_out0), .out1(cmp137_out1));
cmp cmp138 (.in0(cmp138_in0), .in1(cmp138_in1), .out0(cmp138_out0), .out1(cmp138_out1));
cmp cmp139 (.in0(cmp139_in0), .in1(cmp139_in1), .out0(cmp139_out0), .out1(cmp139_out1));
cmp cmp140 (.in0(cmp140_in0), .in1(cmp140_in1), .out0(cmp140_out0), .out1(cmp140_out1));
cmp cmp141 (.in0(cmp141_in0), .in1(cmp141_in1), .out0(cmp141_out0), .out1(cmp141_out1));
cmp cmp142 (.in0(cmp142_in0), .in1(cmp142_in1), .out0(cmp142_out0), .out1(cmp142_out1));
cmp cmp143 (.in0(cmp143_in0), .in1(cmp143_in1), .out0(cmp143_out0), .out1(cmp143_out1));
cmp cmp144 (.in0(cmp144_in0), .in1(cmp144_in1), .out0(cmp144_out0), .out1(cmp144_out1));
cmp cmp145 (.in0(cmp145_in0), .in1(cmp145_in1), .out0(cmp145_out0), .out1(cmp145_out1));
cmp cmp146 (.in0(cmp146_in0), .in1(cmp146_in1), .out0(cmp146_out0), .out1(cmp146_out1));
cmp cmp147 (.in0(cmp147_in0), .in1(cmp147_in1), .out0(cmp147_out0), .out1(cmp147_out1));
cmp cmp148 (.in0(cmp148_in0), .in1(cmp148_in1), .out0(cmp148_out0), .out1(cmp148_out1));
cmp cmp149 (.in0(cmp149_in0), .in1(cmp149_in1), .out0(cmp149_out0), .out1(cmp149_out1));
cmp cmp150 (.in0(cmp150_in0), .in1(cmp150_in1), .out0(cmp150_out0), .out1(cmp150_out1));
cmp cmp151 (.in0(cmp151_in0), .in1(cmp151_in1), .out0(cmp151_out0), .out1(cmp151_out1));
cmp cmp152 (.in0(cmp152_in0), .in1(cmp152_in1), .out0(cmp152_out0), .out1(cmp152_out1));
cmp cmp153 (.in0(cmp153_in0), .in1(cmp153_in1), .out0(cmp153_out0), .out1(cmp153_out1));
cmp cmp154 (.in0(cmp154_in0), .in1(cmp154_in1), .out0(cmp154_out0), .out1(cmp154_out1));
cmp cmp155 (.in0(cmp155_in0), .in1(cmp155_in1), .out0(cmp155_out0), .out1(cmp155_out1));
cmp cmp156 (.in0(cmp156_in0), .in1(cmp156_in1), .out0(cmp156_out0), .out1(cmp156_out1));
cmp cmp157 (.in0(cmp157_in0), .in1(cmp157_in1), .out0(cmp157_out0), .out1(cmp157_out1));
cmp cmp158 (.in0(cmp158_in0), .in1(cmp158_in1), .out0(cmp158_out0), .out1(cmp158_out1));
cmp cmp159 (.in0(cmp159_in0), .in1(cmp159_in1), .out0(cmp159_out0), .out1(cmp159_out1));
cmp cmp160 (.in0(cmp160_in0), .in1(cmp160_in1), .out0(cmp160_out0), .out1(cmp160_out1));
cmp cmp161 (.in0(cmp161_in0), .in1(cmp161_in1), .out0(cmp161_out0), .out1(cmp161_out1));
cmp cmp162 (.in0(cmp162_in0), .in1(cmp162_in1), .out0(cmp162_out0), .out1(cmp162_out1));
cmp cmp163 (.in0(cmp163_in0), .in1(cmp163_in1), .out0(cmp163_out0), .out1(cmp163_out1));
cmp cmp164 (.in0(cmp164_in0), .in1(cmp164_in1), .out0(cmp164_out0), .out1(cmp164_out1));
cmp cmp165 (.in0(cmp165_in0), .in1(cmp165_in1), .out0(cmp165_out0), .out1(cmp165_out1));
cmp cmp166 (.in0(cmp166_in0), .in1(cmp166_in1), .out0(cmp166_out0), .out1(cmp166_out1));
cmp cmp167 (.in0(cmp167_in0), .in1(cmp167_in1), .out0(cmp167_out0), .out1(cmp167_out1));
cmp cmp168 (.in0(cmp168_in0), .in1(cmp168_in1), .out0(cmp168_out0), .out1(cmp168_out1));
cmp cmp169 (.in0(cmp169_in0), .in1(cmp169_in1), .out0(cmp169_out0), .out1(cmp169_out1));
cmp cmp170 (.in0(cmp170_in0), .in1(cmp170_in1), .out0(cmp170_out0), .out1(cmp170_out1));
cmp cmp171 (.in0(cmp171_in0), .in1(cmp171_in1), .out0(cmp171_out0), .out1(cmp171_out1));
cmp cmp172 (.in0(cmp172_in0), .in1(cmp172_in1), .out0(cmp172_out0), .out1(cmp172_out1));
cmp cmp173 (.in0(cmp173_in0), .in1(cmp173_in1), .out0(cmp173_out0), .out1(cmp173_out1));
cmp cmp174 (.in0(cmp174_in0), .in1(cmp174_in1), .out0(cmp174_out0), .out1(cmp174_out1));
cmp cmp175 (.in0(cmp175_in0), .in1(cmp175_in1), .out0(cmp175_out0), .out1(cmp175_out1));
cmp cmp176 (.in0(cmp176_in0), .in1(cmp176_in1), .out0(cmp176_out0), .out1(cmp176_out1));
cmp cmp177 (.in0(cmp177_in0), .in1(cmp177_in1), .out0(cmp177_out0), .out1(cmp177_out1));
cmp cmp178 (.in0(cmp178_in0), .in1(cmp178_in1), .out0(cmp178_out0), .out1(cmp178_out1));
cmp cmp179 (.in0(cmp179_in0), .in1(cmp179_in1), .out0(cmp179_out0), .out1(cmp179_out1));
cmp cmp180 (.in0(cmp180_in0), .in1(cmp180_in1), .out0(cmp180_out0), .out1(cmp180_out1));
cmp cmp181 (.in0(cmp181_in0), .in1(cmp181_in1), .out0(cmp181_out0), .out1(cmp181_out1));
cmp cmp182 (.in0(cmp182_in0), .in1(cmp182_in1), .out0(cmp182_out0), .out1(cmp182_out1));
cmp cmp183 (.in0(cmp183_in0), .in1(cmp183_in1), .out0(cmp183_out0), .out1(cmp183_out1));
cmp cmp184 (.in0(cmp184_in0), .in1(cmp184_in1), .out0(cmp184_out0), .out1(cmp184_out1));
cmp cmp185 (.in0(cmp185_in0), .in1(cmp185_in1), .out0(cmp185_out0), .out1(cmp185_out1));
cmp cmp186 (.in0(cmp186_in0), .in1(cmp186_in1), .out0(cmp186_out0), .out1(cmp186_out1));
cmp cmp187 (.in0(cmp187_in0), .in1(cmp187_in1), .out0(cmp187_out0), .out1(cmp187_out1));
cmp cmp188 (.in0(cmp188_in0), .in1(cmp188_in1), .out0(cmp188_out0), .out1(cmp188_out1));
cmp cmp189 (.in0(cmp189_in0), .in1(cmp189_in1), .out0(cmp189_out0), .out1(cmp189_out1));
cmp cmp190 (.in0(cmp190_in0), .in1(cmp190_in1), .out0(cmp190_out0), .out1(cmp190_out1));
cmp cmp191 (.in0(cmp191_in0), .in1(cmp191_in1), .out0(cmp191_out0), .out1(cmp191_out1));
cmp cmp192 (.in0(cmp192_in0), .in1(cmp192_in1), .out0(cmp192_out0), .out1(cmp192_out1));
cmp cmp193 (.in0(cmp193_in0), .in1(cmp193_in1), .out0(cmp193_out0), .out1(cmp193_out1));
cmp cmp194 (.in0(cmp194_in0), .in1(cmp194_in1), .out0(cmp194_out0), .out1(cmp194_out1));
cmp cmp195 (.in0(cmp195_in0), .in1(cmp195_in1), .out0(cmp195_out0), .out1(cmp195_out1));
cmp cmp196 (.in0(cmp196_in0), .in1(cmp196_in1), .out0(cmp196_out0), .out1(cmp196_out1));
cmp cmp197 (.in0(cmp197_in0), .in1(cmp197_in1), .out0(cmp197_out0), .out1(cmp197_out1));
cmp cmp198 (.in0(cmp198_in0), .in1(cmp198_in1), .out0(cmp198_out0), .out1(cmp198_out1));
cmp cmp199 (.in0(cmp199_in0), .in1(cmp199_in1), .out0(cmp199_out0), .out1(cmp199_out1));
cmp cmp200 (.in0(cmp200_in0), .in1(cmp200_in1), .out0(cmp200_out0), .out1(cmp200_out1));
cmp cmp201 (.in0(cmp201_in0), .in1(cmp201_in1), .out0(cmp201_out0), .out1(cmp201_out1));
cmp cmp202 (.in0(cmp202_in0), .in1(cmp202_in1), .out0(cmp202_out0), .out1(cmp202_out1));
cmp cmp203 (.in0(cmp203_in0), .in1(cmp203_in1), .out0(cmp203_out0), .out1(cmp203_out1));
cmp cmp204 (.in0(cmp204_in0), .in1(cmp204_in1), .out0(cmp204_out0), .out1(cmp204_out1));
cmp cmp205 (.in0(cmp205_in0), .in1(cmp205_in1), .out0(cmp205_out0), .out1(cmp205_out1));
cmp cmp206 (.in0(cmp206_in0), .in1(cmp206_in1), .out0(cmp206_out0), .out1(cmp206_out1));
cmp cmp207 (.in0(cmp207_in0), .in1(cmp207_in1), .out0(cmp207_out0), .out1(cmp207_out1));
cmp cmp208 (.in0(cmp208_in0), .in1(cmp208_in1), .out0(cmp208_out0), .out1(cmp208_out1));
cmp cmp209 (.in0(cmp209_in0), .in1(cmp209_in1), .out0(cmp209_out0), .out1(cmp209_out1));
cmp cmp210 (.in0(cmp210_in0), .in1(cmp210_in1), .out0(cmp210_out0), .out1(cmp210_out1));
cmp cmp211 (.in0(cmp211_in0), .in1(cmp211_in1), .out0(cmp211_out0), .out1(cmp211_out1));
cmp cmp212 (.in0(cmp212_in0), .in1(cmp212_in1), .out0(cmp212_out0), .out1(cmp212_out1));
cmp cmp213 (.in0(cmp213_in0), .in1(cmp213_in1), .out0(cmp213_out0), .out1(cmp213_out1));
cmp cmp214 (.in0(cmp214_in0), .in1(cmp214_in1), .out0(cmp214_out0), .out1(cmp214_out1));
cmp cmp215 (.in0(cmp215_in0), .in1(cmp215_in1), .out0(cmp215_out0), .out1(cmp215_out1));
cmp cmp216 (.in0(cmp216_in0), .in1(cmp216_in1), .out0(cmp216_out0), .out1(cmp216_out1));
cmp cmp217 (.in0(cmp217_in0), .in1(cmp217_in1), .out0(cmp217_out0), .out1(cmp217_out1));
cmp cmp218 (.in0(cmp218_in0), .in1(cmp218_in1), .out0(cmp218_out0), .out1(cmp218_out1));
cmp cmp219 (.in0(cmp219_in0), .in1(cmp219_in1), .out0(cmp219_out0), .out1(cmp219_out1));
cmp cmp220 (.in0(cmp220_in0), .in1(cmp220_in1), .out0(cmp220_out0), .out1(cmp220_out1));
cmp cmp221 (.in0(cmp221_in0), .in1(cmp221_in1), .out0(cmp221_out0), .out1(cmp221_out1));
cmp cmp222 (.in0(cmp222_in0), .in1(cmp222_in1), .out0(cmp222_out0), .out1(cmp222_out1));
cmp cmp223 (.in0(cmp223_in0), .in1(cmp223_in1), .out0(cmp223_out0), .out1(cmp223_out1));
cmp cmp224 (.in0(cmp224_in0), .in1(cmp224_in1), .out0(cmp224_out0), .out1(cmp224_out1));
cmp cmp225 (.in0(cmp225_in0), .in1(cmp225_in1), .out0(cmp225_out0), .out1(cmp225_out1));
cmp cmp226 (.in0(cmp226_in0), .in1(cmp226_in1), .out0(cmp226_out0), .out1(cmp226_out1));
cmp cmp227 (.in0(cmp227_in0), .in1(cmp227_in1), .out0(cmp227_out0), .out1(cmp227_out1));
cmp cmp228 (.in0(cmp228_in0), .in1(cmp228_in1), .out0(cmp228_out0), .out1(cmp228_out1));
cmp cmp229 (.in0(cmp229_in0), .in1(cmp229_in1), .out0(cmp229_out0), .out1(cmp229_out1));
cmp cmp230 (.in0(cmp230_in0), .in1(cmp230_in1), .out0(cmp230_out0), .out1(cmp230_out1));
cmp cmp231 (.in0(cmp231_in0), .in1(cmp231_in1), .out0(cmp231_out0), .out1(cmp231_out1));
cmp cmp232 (.in0(cmp232_in0), .in1(cmp232_in1), .out0(cmp232_out0), .out1(cmp232_out1));
cmp cmp233 (.in0(cmp233_in0), .in1(cmp233_in1), .out0(cmp233_out0), .out1(cmp233_out1));
cmp cmp234 (.in0(cmp234_in0), .in1(cmp234_in1), .out0(cmp234_out0), .out1(cmp234_out1));
cmp cmp235 (.in0(cmp235_in0), .in1(cmp235_in1), .out0(cmp235_out0), .out1(cmp235_out1));
cmp cmp236 (.in0(cmp236_in0), .in1(cmp236_in1), .out0(cmp236_out0), .out1(cmp236_out1));
cmp cmp237 (.in0(cmp237_in0), .in1(cmp237_in1), .out0(cmp237_out0), .out1(cmp237_out1));
cmp cmp238 (.in0(cmp238_in0), .in1(cmp238_in1), .out0(cmp238_out0), .out1(cmp238_out1));
cmp cmp239 (.in0(cmp239_in0), .in1(cmp239_in1), .out0(cmp239_out0), .out1(cmp239_out1));
cmp cmp240 (.in0(cmp240_in0), .in1(cmp240_in1), .out0(cmp240_out0), .out1(cmp240_out1));
cmp cmp241 (.in0(cmp241_in0), .in1(cmp241_in1), .out0(cmp241_out0), .out1(cmp241_out1));
cmp cmp242 (.in0(cmp242_in0), .in1(cmp242_in1), .out0(cmp242_out0), .out1(cmp242_out1));
cmp cmp243 (.in0(cmp243_in0), .in1(cmp243_in1), .out0(cmp243_out0), .out1(cmp243_out1));
cmp cmp244 (.in0(cmp244_in0), .in1(cmp244_in1), .out0(cmp244_out0), .out1(cmp244_out1));
cmp cmp245 (.in0(cmp245_in0), .in1(cmp245_in1), .out0(cmp245_out0), .out1(cmp245_out1));
cmp cmp246 (.in0(cmp246_in0), .in1(cmp246_in1), .out0(cmp246_out0), .out1(cmp246_out1));
cmp cmp247 (.in0(cmp247_in0), .in1(cmp247_in1), .out0(cmp247_out0), .out1(cmp247_out1));
cmp cmp248 (.in0(cmp248_in0), .in1(cmp248_in1), .out0(cmp248_out0), .out1(cmp248_out1));
cmp cmp249 (.in0(cmp249_in0), .in1(cmp249_in1), .out0(cmp249_out0), .out1(cmp249_out1));
cmp cmp250 (.in0(cmp250_in0), .in1(cmp250_in1), .out0(cmp250_out0), .out1(cmp250_out1));
cmp cmp251 (.in0(cmp251_in0), .in1(cmp251_in1), .out0(cmp251_out0), .out1(cmp251_out1));
cmp cmp252 (.in0(cmp252_in0), .in1(cmp252_in1), .out0(cmp252_out0), .out1(cmp252_out1));
cmp cmp253 (.in0(cmp253_in0), .in1(cmp253_in1), .out0(cmp253_out0), .out1(cmp253_out1));
cmp cmp254 (.in0(cmp254_in0), .in1(cmp254_in1), .out0(cmp254_out0), .out1(cmp254_out1));
cmp cmp255 (.in0(cmp255_in0), .in1(cmp255_in1), .out0(cmp255_out0), .out1(cmp255_out1));
cmp cmp256 (.in0(cmp256_in0), .in1(cmp256_in1), .out0(cmp256_out0), .out1(cmp256_out1));
cmp cmp257 (.in0(cmp257_in0), .in1(cmp257_in1), .out0(cmp257_out0), .out1(cmp257_out1));
cmp cmp258 (.in0(cmp258_in0), .in1(cmp258_in1), .out0(cmp258_out0), .out1(cmp258_out1));
cmp cmp259 (.in0(cmp259_in0), .in1(cmp259_in1), .out0(cmp259_out0), .out1(cmp259_out1));
cmp cmp260 (.in0(cmp260_in0), .in1(cmp260_in1), .out0(cmp260_out0), .out1(cmp260_out1));
cmp cmp261 (.in0(cmp261_in0), .in1(cmp261_in1), .out0(cmp261_out0), .out1(cmp261_out1));
cmp cmp262 (.in0(cmp262_in0), .in1(cmp262_in1), .out0(cmp262_out0), .out1(cmp262_out1));
cmp cmp263 (.in0(cmp263_in0), .in1(cmp263_in1), .out0(cmp263_out0), .out1(cmp263_out1));
cmp cmp264 (.in0(cmp264_in0), .in1(cmp264_in1), .out0(cmp264_out0), .out1(cmp264_out1));
cmp cmp265 (.in0(cmp265_in0), .in1(cmp265_in1), .out0(cmp265_out0), .out1(cmp265_out1));
cmp cmp266 (.in0(cmp266_in0), .in1(cmp266_in1), .out0(cmp266_out0), .out1(cmp266_out1));
cmp cmp267 (.in0(cmp267_in0), .in1(cmp267_in1), .out0(cmp267_out0), .out1(cmp267_out1));
cmp cmp268 (.in0(cmp268_in0), .in1(cmp268_in1), .out0(cmp268_out0), .out1(cmp268_out1));
cmp cmp269 (.in0(cmp269_in0), .in1(cmp269_in1), .out0(cmp269_out0), .out1(cmp269_out1));
cmp cmp270 (.in0(cmp270_in0), .in1(cmp270_in1), .out0(cmp270_out0), .out1(cmp270_out1));
cmp cmp271 (.in0(cmp271_in0), .in1(cmp271_in1), .out0(cmp271_out0), .out1(cmp271_out1));
cmp cmp272 (.in0(cmp272_in0), .in1(cmp272_in1), .out0(cmp272_out0), .out1(cmp272_out1));
cmp cmp273 (.in0(cmp273_in0), .in1(cmp273_in1), .out0(cmp273_out0), .out1(cmp273_out1));
cmp cmp274 (.in0(cmp274_in0), .in1(cmp274_in1), .out0(cmp274_out0), .out1(cmp274_out1));
cmp cmp275 (.in0(cmp275_in0), .in1(cmp275_in1), .out0(cmp275_out0), .out1(cmp275_out1));
cmp cmp276 (.in0(cmp276_in0), .in1(cmp276_in1), .out0(cmp276_out0), .out1(cmp276_out1));
cmp cmp277 (.in0(cmp277_in0), .in1(cmp277_in1), .out0(cmp277_out0), .out1(cmp277_out1));
cmp cmp278 (.in0(cmp278_in0), .in1(cmp278_in1), .out0(cmp278_out0), .out1(cmp278_out1));
cmp cmp279 (.in0(cmp279_in0), .in1(cmp279_in1), .out0(cmp279_out0), .out1(cmp279_out1));
cmp cmp280 (.in0(cmp280_in0), .in1(cmp280_in1), .out0(cmp280_out0), .out1(cmp280_out1));
cmp cmp281 (.in0(cmp281_in0), .in1(cmp281_in1), .out0(cmp281_out0), .out1(cmp281_out1));
cmp cmp282 (.in0(cmp282_in0), .in1(cmp282_in1), .out0(cmp282_out0), .out1(cmp282_out1));
cmp cmp283 (.in0(cmp283_in0), .in1(cmp283_in1), .out0(cmp283_out0), .out1(cmp283_out1));
cmp cmp284 (.in0(cmp284_in0), .in1(cmp284_in1), .out0(cmp284_out0), .out1(cmp284_out1));
cmp cmp285 (.in0(cmp285_in0), .in1(cmp285_in1), .out0(cmp285_out0), .out1(cmp285_out1));
cmp cmp286 (.in0(cmp286_in0), .in1(cmp286_in1), .out0(cmp286_out0), .out1(cmp286_out1));
cmp cmp287 (.in0(cmp287_in0), .in1(cmp287_in1), .out0(cmp287_out0), .out1(cmp287_out1));
cmp cmp288 (.in0(cmp288_in0), .in1(cmp288_in1), .out0(cmp288_out0), .out1(cmp288_out1));
cmp cmp289 (.in0(cmp289_in0), .in1(cmp289_in1), .out0(cmp289_out0), .out1(cmp289_out1));
cmp cmp290 (.in0(cmp290_in0), .in1(cmp290_in1), .out0(cmp290_out0), .out1(cmp290_out1));
cmp cmp291 (.in0(cmp291_in0), .in1(cmp291_in1), .out0(cmp291_out0), .out1(cmp291_out1));
cmp cmp292 (.in0(cmp292_in0), .in1(cmp292_in1), .out0(cmp292_out0), .out1(cmp292_out1));
cmp cmp293 (.in0(cmp293_in0), .in1(cmp293_in1), .out0(cmp293_out0), .out1(cmp293_out1));
cmp cmp294 (.in0(cmp294_in0), .in1(cmp294_in1), .out0(cmp294_out0), .out1(cmp294_out1));
cmp cmp295 (.in0(cmp295_in0), .in1(cmp295_in1), .out0(cmp295_out0), .out1(cmp295_out1));
cmp cmp296 (.in0(cmp296_in0), .in1(cmp296_in1), .out0(cmp296_out0), .out1(cmp296_out1));
cmp cmp297 (.in0(cmp297_in0), .in1(cmp297_in1), .out0(cmp297_out0), .out1(cmp297_out1));
cmp cmp298 (.in0(cmp298_in0), .in1(cmp298_in1), .out0(cmp298_out0), .out1(cmp298_out1));
cmp cmp299 (.in0(cmp299_in0), .in1(cmp299_in1), .out0(cmp299_out0), .out1(cmp299_out1));
cmp cmp300 (.in0(cmp300_in0), .in1(cmp300_in1), .out0(cmp300_out0), .out1(cmp300_out1));
cmp cmp301 (.in0(cmp301_in0), .in1(cmp301_in1), .out0(cmp301_out0), .out1(cmp301_out1));
cmp cmp302 (.in0(cmp302_in0), .in1(cmp302_in1), .out0(cmp302_out0), .out1(cmp302_out1));
cmp cmp303 (.in0(cmp303_in0), .in1(cmp303_in1), .out0(cmp303_out0), .out1(cmp303_out1));
cmp cmp304 (.in0(cmp304_in0), .in1(cmp304_in1), .out0(cmp304_out0), .out1(cmp304_out1));
cmp cmp305 (.in0(cmp305_in0), .in1(cmp305_in1), .out0(cmp305_out0), .out1(cmp305_out1));
cmp cmp306 (.in0(cmp306_in0), .in1(cmp306_in1), .out0(cmp306_out0), .out1(cmp306_out1));
cmp cmp307 (.in0(cmp307_in0), .in1(cmp307_in1), .out0(cmp307_out0), .out1(cmp307_out1));
cmp cmp308 (.in0(cmp308_in0), .in1(cmp308_in1), .out0(cmp308_out0), .out1(cmp308_out1));
cmp cmp309 (.in0(cmp309_in0), .in1(cmp309_in1), .out0(cmp309_out0), .out1(cmp309_out1));
cmp cmp310 (.in0(cmp310_in0), .in1(cmp310_in1), .out0(cmp310_out0), .out1(cmp310_out1));
cmp cmp311 (.in0(cmp311_in0), .in1(cmp311_in1), .out0(cmp311_out0), .out1(cmp311_out1));
cmp cmp312 (.in0(cmp312_in0), .in1(cmp312_in1), .out0(cmp312_out0), .out1(cmp312_out1));
endmodule

module cmp(
     input  [7:0] in0,
     input  [7:0] in1,
     output wire [7:0] out0,
     output wire [7:0] out1
);
     assign out0 = (in0<in1) ? in0:in1;
     assign out1 = (in0<in1) ? in1:in0;
endmodule
